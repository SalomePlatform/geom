-- Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	NMTTools_CommonBlockAPI.cdl
-- Created:	Mon Dec 15 11:35:46 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class CommonBlockAPI from NMTTools 

	---Purpose: 

uses
    ListOfCommonBlock from NMTTools, 
    ListOfPaveBlock   from BOPTools, 
    PaveBlock         from BOPTools, 
    CommonBlock       from NMTTools 
    
--raises

is 
    Create  (aList:ListOfCommonBlock from NMTTools)   
    	returns CommonBlockAPI from NMTTools; 
	 
    List(me) 
    	returns  ListOfCommonBlock from NMTTools; 
    ---C++:  return const & 
    	---Purpose:   
    	--- Selector 
    	---
    CommonPaveBlocks(me;   
    	    anE:Integer from  Standard) 
    	returns  ListOfPaveBlock from BOPTools;
    ---C++:  return const &  
    	---Purpose:   
    	--- Returns all PaveBlock-s (from the list) that are 
    	--- common for the given edge with  DS-index <anE>     
    	---
    IsCommonBlock   (me;  
    	    aPB: PaveBlock from BOPTools) 
    	returns  Boolean from Standard;
    	---Purpose:   
    	--- Returns TRUE if given PaveBlock <aPB> is 
    	--- common for the Blocks from the list  
	 
    CommonBlock(me; 
    	    aPB: PaveBlock from BOPTools) 
	returns  CommonBlock from NMTTools;  
    ---C++:  return &     

fields
    myListOfCommonBlock  :Address from Standard;
    myListOfPaveBlock    :ListOfPaveBlock from BOPTools;
    
end CommonBlockAPI;
