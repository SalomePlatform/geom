-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	GEOMAlgo_ShapeInfo.cdl
--  Created:	Mon Apr  2 14:04:24 2007
--  Author:	Peter KURNEV
--
class ShapeInfo from GEOMAlgo 

	---Purpose: 

uses 
    Pnt from gp, 
    Dir from gp, 
    Ax2 from gp, 
    Ax3 from gp, 
    
    ShapeEnum from TopAbs, 
    Shape from TopoDS, 
     
    KindOfShape   from GEOMAlgo,
    KindOfBounds  from GEOMAlgo, 
    KindOfClosed  from GEOMAlgo, 
    KindOfName from GEOMAlgo
--raises

is 
    Create 
    	returns ShapeInfo from GEOMAlgo;   
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_ShapeInfo();" 
     
    Reset(me:out); 
     
    SetType(me:out; 
    	    aType:ShapeEnum from TopAbs); 
	 
    Type(me) 
    	returns ShapeEnum from TopAbs; 
	 
    SetNbSubShapes(me:out; 
    	    aType:ShapeEnum from TopAbs; 
    	    aNb  :Integer from Standard); 
     
    NbSubShapes(me; 
    	    aType:ShapeEnum from TopAbs) 
    	returns Integer from Standard; 
	 
    SetKindOfShape (me:out; 
    	    aT:KindOfShape from GEOMAlgo); 
	 
    KindOfShape (me) 
    	 returns KindOfShape from GEOMAlgo;      

    SetKindOfName (me:out; 
    	    aT: KindOfName from GEOMAlgo); 
	 
    KindOfName(me) 
    	 returns KindOfName from GEOMAlgo; 

    SetKindOfBounds (me:out; 
    	    aT:KindOfBounds from GEOMAlgo); 
	     
    KindOfBounds (me) 
    	 returns KindOfBounds from GEOMAlgo;    
	  
    SetKindOfClosed (me:out; 
    	    aT:KindOfClosed from GEOMAlgo); 
	     
    KindOfClosed(me) 
    	 returns KindOfClosed from GEOMAlgo;   
	 
    SetLocation (me:out; 
    	    aP: Pnt from gp); 
	     
    Location (me) 
    	 returns Pnt from gp; 
    ---C++: return const&  
	 
    SetDirection  (me:out; 
    	    aD:Dir from gp); 
	     
    Direction  (me) 
    	 returns Dir from gp; 
    ---C++: return const&      
      
    SetPosition (me:out;  
    	    aAx2 : Ax2 from gp);
     
    SetPosition (me:out;  
    	    aAx3 : Ax3 from gp); 
	 
    Position (me)  
    	returns Ax3 from gp; 
    ---C++: return const&	   
  	
    SetPnt1 (me:out; 
    	    aP: Pnt from gp); 
	     
    Pnt1 (me) 
    	 returns Pnt from gp; 
    ---C++: return const& 
     
    SetPnt2 (me:out; 
    	    aP: Pnt from gp); 
	     
    Pnt2 (me) 
    	 returns Pnt from gp; 
    ---C++: return const& 
     
    SetRadius1 (me:out; 
    	    aR: Real from Standard); 
	     
    Radius1(me) 
    	 returns Real from Standard;    

    SetRadius2 (me:out; 
    	    aR: Real from Standard); 
	     
    Radius2(me) 
    	 returns Real from Standard;   
      
    SetLength(me:out; 
    	    aL: Real from Standard); 
	     
    Length(me) 
    	 returns Real from Standard;  
	  
    SetWidth(me:out; 
    	    aW: Real from Standard); 
	     
    Width(me) 
    	 returns Real from Standard;  
	   
    SetHeight(me:out; 
    	    aH: Real from Standard); 
	     
    Height(me) 
    	 returns Real from Standard; 
    --
    -- Dump
    --  	     
    Dump(me); 
    	
    DumpVertex(me) 
    	is protected; 
	 
    DumpEdge(me) 
    	is protected; 
	 
    DumpWire(me) 
    	is protected;
  
    DumpFace(me) 
    	is protected;
  
    DumpShell(me) 
    	is protected; 
     
    DumpSolid(me) 
    	is protected; 
	 
    DumpCompSolid(me) 
    	is protected; 
	 
    DumpCompound(me) 
    	is protected;
 
fields 
    myType          : ShapeEnum from TopAbs      is protected; 
    myNbSubShapes   : Integer from Standard[9]   is protected; 
    myKindOfShape   : KindOfShape from GEOMAlgo  is protected;  
    myKindOfName    : KindOfName from GEOMAlgo   is protected;  
    myKindOfBounds  : KindOfBounds from GEOMAlgo is protected;  
    myKindOfClosed  : KindOfClosed from GEOMAlgo is protected;  
    --
    myLocation      : Pnt from gp is protected;  
    myDirection     : Dir from gp is protected; 
    myPosition      : Ax3 from gp is protected; 
    -- 
    myRadius1       : Real from Standard is protected;    
    myRadius2       : Real from Standard is protected;    
    myLength        : Real from Standard is protected;    
    myWidth         : Real from Standard is protected;    
    myHeight        : Real from Standard is protected;    
    -- 
    myPnt1          : Pnt from gp is protected;   
    myPnt2          : Pnt from gp is protected;    
    -- 
    myNbTypes       : Integer from Standard is protected;
end ShapeInfo;
