--  Copyright (C) 2007-2010  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	NMTDS_PassKeyBoolean.cdl
--  Created:	
--  Author:	Peter KURNEV
--
class PassKeyBoolean from NMTDS 
    inherits  PassKey from NMTDS 

	---Purpose: 

uses
    Shape from TopoDS, 
    ListOfInteger from TColStd   
  	 
--raises

is 
    Create  
    	returns PassKeyBoolean from NMTDS; 
    ---C++: alias "Standard_EXPORT virtual ~NMTDS_PassKeyBoolean();" 
    
    SetFlag(me:out; 
    	    aFlag: Boolean from Standard); 
    ---C++: alias " Standard_EXPORT NMTDS_PassKeyBoolean& operator =(const NMTDS_PassKeyBoolean& Other);" 
    
    Flag(me)  
    	returns Boolean from Standard;      

fields 
    myFlag: Boolean from Standard is protected;  

end PassKeyBoolean;
