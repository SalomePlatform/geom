// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
// See http://www.salome-platform.org/
//
-- File:	NMTTools_PCurveMaker.cdl
-- Created:	 
-- Author:	Peter KURNEV
--		<pkv@irinox>

class PCurveMaker from NMTTools 

	---Purpose:  
    	--  Class provides computation p-curves for the edges and theirs  
        --- split parts  	

uses 
    PDSFiller from NMTTools
    
is   
    Create (aFiller:out PDSFiller from NMTTools)  
    	returns PCurveMaker from NMTTools; 
    	---Purpose:  
    	--- Constructor 
    	---
    Do(me:out);   
    	---Purpose: 
    	--- Launch the processor   
    	---
    IsDone(me) 
    	returns Boolean from Standard;  
    	---Purpose:  
    	--- Returns TRUE if Ok       
    	---
	
fields  
    myDSFiller: PDSFiller from NMTTools  	is protected;
    myIsDone  : Boolean   from Standard	        is protected;   
    
end PCurveMaker;
