// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
// See http://www.salome-platform.org/
//
-- File:	NMTAlgo.cdl
-- Created:	Tue Jan 27 14:39:05 2004
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2004


package NMTAlgo 

	---Purpose: 

uses
    TCollection,
    TColStd, 
    gp,
    TopAbs, 
    TopoDS, 
    TopTools,  
    
    BooleanOperations,
    BOPTColStd,
    IntTools,
    BOPTools, 
    BOP, 
     
    NMTDS,
    NMTTools, 
      
    BRep,
    BRepAlgo 
    
is 
    deferred class Algo; 
    class Splitter; 
    class Splitter1; --modified by NIZNHY-PKV Wed Feb 11 14:28:50 2004
    class Builder; 
    class Tools; 
    class Loop3d; 
      	
end NMTAlgo;
