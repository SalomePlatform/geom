-- Copyright (C) 2007-2019  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License, or (at your option) any later version.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
-- File:	GEOMAlgo.cdl
-- Created:	Sat Dec 04 12:36:22 2004
-- Author:	Peter KURNEV

package GEOMAlgo

	---Purpose:

--uses
 
is
    --  Enumerations
    imported State from GEOMAlgo;
    imported KindOfShape from GEOMAlgo;
    imported KindOfName from GEOMAlgo;
    imported KindOfBounds from GEOMAlgo;
    imported KindOfClosed from GEOMAlgo;
    --  
    -- Algos 
    -- 
    imported Algo from GEOMAlgo;
    imported ShapeSolid from GEOMAlgo;  
    imported VertexSolid from GEOMAlgo;  
    imported WireSolid from GEOMAlgo; 
    imported ShellSolid from GEOMAlgo; 
    imported SolidSolid from GEOMAlgo;  
    imported FinderShapeOn from GEOMAlgo; 
    imported FinderShapeOn1 from GEOMAlgo; 
    imported HAlgo from GEOMAlgo; 
    imported ShapeAlgo from GEOMAlgo;  
    imported Clsf from GEOMAlgo; 
    imported ClsfBox from GEOMAlgo;  
    imported ClsfSurf from GEOMAlgo;
    imported ClsfSolid from GEOMAlgo; 
    imported FinderShapeOn2 from GEOMAlgo;
    imported FinderShapeOnQuad from GEOMAlgo; 
    imported Gluer from GEOMAlgo; 
    imported GlueAnalyser from GEOMAlgo; 
    imported GluerAlgo from GEOMAlgo; 
    imported GlueDetector from GEOMAlgo; 
    imported BuilderShape from GEOMAlgo;
    imported Gluer2 from GEOMAlgo; 
    imported GetInPlace from GEOMAlgo; 
    imported Splitter from GEOMAlgo;
    --  
    
    -- 
    imported AlgoTools from GEOMAlgo;
     
    --  Gluer / GetInPlace
    --
    
    
    --
    -- Algos
    imported RemoverWebs from GEOMAlgo;

    --imported WireSplitter from GEOMAlgo;
    --imported WESScaler from GEOMAlgo;
    --imported WESCorrector from GEOMAlgo;
    --imported WireEdgeSet from GEOMAlgo;
    --imported GlueAnalyser from GEOMAlgo;
    --imported Gluer from GEOMAlgo;
    
    --
    
    --imported Splitter from GEOMAlgo;
    --imported Builder from GEOMAlgo;
    
    --imported BuilderSolid from GEOMAlgo;
    --imported BuilderFace from GEOMAlgo;
    --imported BuilderArea from GEOMAlgo;

    imported ShapeInfoFiller from GEOMAlgo;
    --
    -- Data /  Tools
    --imported ShapeSet from GEOMAlgo;
    imported SurfaceTools from GEOMAlgo;
    imported ShapeInfo from GEOMAlgo;
    imported CoupleOfShapes from GEOMAlgo;
    --imported BuilderTools from GEOMAlgo;
    --imported Tools3D from GEOMAlgo;
    --imported Tools from GEOMAlgo;
    --imported PWireEdgeSet from GEOMAlgo;
    imported BndSphere from GEOMAlgo;
    imported StateCollector from GEOMAlgo;
    imported PassKey from GEOMAlgo;
    imported PassKeyMapHasher from GEOMAlgo;
    imported PassKeyShape from GEOMAlgo;
    imported PassKeyShapeMapHasher from GEOMAlgo;
    imported ListOfCoupleOfShapes from GEOMAlgo;
    imported ListIteratorOfListOfCoupleOfShapes from GEOMAlgo;
    imported ListOfPnt from GEOMAlgo;
    imported ListIteratorOfListOfPnt from GEOMAlgo; 
    imported IndexedDataMapOfShapeIndexedMapOfShape from GEOMAlgo; 
    
    --imported DataMapOfShapeShapeSet from GEOMAlgo;
    --imported DataMapIteratorOfDataMapOfShapeShapeSet from GEOMAlgo;
    --imported DataMapOfShapeReal from GEOMAlgo;
    --imported DataMapIteratorOfDataMapOfShapeReal from GEOMAlgo;
    --imported DataMapOfRealListOfShape from GEOMAlgo;
    --imported DataMapIteratorOfDataMapOfRealListOfShape from GEOMAlgo;
    imported DataMapOfPassKeyInteger from GEOMAlgo;
    imported DataMapIteratorOfDataMapOfPassKeyInteger from GEOMAlgo;
    --imported DataMapOfPassKeyShapeShape from GEOMAlgo;
    --imported DataMapIteratorOfDataMapOfPassKeyShapeShape from GEOMAlgo;
    --imported DataMapOfOrientedShapeShape from GEOMAlgo;
    --imported DataMapIteratorOfDataMapOfOrientedShapeShape from GEOMAlgo;
    imported DataMapOfShapeMapOfShape from GEOMAlgo;
    imported DataMapIteratorOfDataMapOfShapeMapOfShape from GEOMAlgo;
    imported DataMapOfShapePnt from GEOMAlgo;
    imported DataMapIteratorOfDataMapOfShapePnt from GEOMAlgo;
    imported IndexedDataMapOfShapeBox from GEOMAlgo;
    imported IndexedDataMapOfShapeShapeInfo from GEOMAlgo;
    imported IndexedDataMapOfShapeState from GEOMAlgo;
    imported IndexedDataMapOfIntegerShape from GEOMAlgo;
    imported IndexedDataMapOfPassKeyShapeListOfShape from GEOMAlgo;

end GEOMAlgo;
