--  Copyright (C) 2007-2010  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	NMTTools_DSFiller.cdl
-- Created:	Fri Dec  5 13:57:03 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class DSFiller from NMTTools 

	---Purpose: 

uses
    Shape from TopoDS,  
    InterferencePool     from BOPTools, 
    PInterferencePool    from BOPTools,
    ShapesDataStructure  from NMTDS, 
    PShapesDataStructure from NMTDS,
    PPaveFiller          from NMTTools, 
    PaveFiller           from NMTTools
--raises

is  
    Create  
    	returns DSFiller from NMTTools; 
	 
    Destroy (me:out);
    ---C++: alias ~
    ---Purpose: Destructor 
    -- 
    --  Selectors/Modifiers   
    SetCompositeShape (me:out;  
    	    aS:  Shape from TopoDS);  
     
    CompositeShape(me) 
    	returns  Shape from TopoDS; 
    	---C++:  return  const& 
     
    SetNewFiller(me;  
    	    aFlag:Boolean from  Standard); 
     
    IsNewFiller(me) 
    	returns Boolean from  Standard;  
    --	 
    --  Perform the algo      
    Perform (me:out);   
    --
    --  Protected section 
    Clear   (me:out) 
    	is protected;  
    --
    -- Query section 
    DS  (me) 
	returns  ShapesDataStructure from NMTDS; 
    	---C++:  return const &    
	 
    InterfPool (me) 
    	returns  InterferencePool from BOPTools;
    ---C++:  return const & 
	 
    IsDone(me) 
    	returns  Boolean  from  Standard; 
      
    PaveFiller(me) 
	returns PaveFiller from NMTTools; 
    ---C++:  return const &

    ChangePaveFiller (me:out) 
	returns PaveFiller from NMTTools; 
    ---C++:  return &

fields
    myCompositeShape  :  Shape from TopoDS is protected;
    myDS              :  PShapesDataStructure from NMTDS is protected; 
    myInterfPool      :  PInterferencePool    from BOPTools is protected;  
    myPaveFiller      :  PPaveFiller from NMTTools is protected;   

    myIsDone          :  Boolean from  Standard is protected; 
    myIsNewFiller     :  Boolean from  Standard is protected;  

end DSFiller;
