-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	NMTDS.cdl
--  Created:	Fri Nov 28 10:13:19 2003
--  Author:	Peter KURNEV
--
package NMTDS 

	---Purpose: 

--uses   
    --TCollection, 
    --TColStd,
    --gp,
    --Bnd,
    --TopoDS, 
    --TopAbs, 
    --TopTools, 
    --BooleanOperations, 
    --BOPTools,
    --BOPTColStd 
    
is  
    imported InterfType from NMTDS; 
    imported BndSphere from NMTDS; 
    imported IndexRange from NMTDS;
    imported InterfPool from NMTDS;
    imported Iterator from NMTDS;
    imported IteratorCheckerSI from NMTDS;
    imported Pair from NMTDS;
    imported PairBoolean from NMTDS;
    imported PairMapHasher from NMTDS;
    imported PassKey from NMTDS;
    imported PassKeyBoolean from NMTDS;
    imported PassKeyMapHasher from NMTDS;
    imported PassKeyShape from NMTDS;
    imported PassKeyShapeMapHasher from NMTDS;
    imported Tools from NMTDS;
    imported ShapesDataStructure from NMTDS;
    imported PShapesDataStructure from NMTDS;
    imported PIterator from NMTDS;
    imported PInterfPool from NMTDS;  
    --
    imported ListOfPassKey from NMTDS;
    imported ListIteratorOfListOfPassKey  from NMTDS;
 
    imported ListOfPassKeyBoolean from NMTDS;
    imported ListIteratorOfListOfPassKeyBoolean from NMTDS;  
     
    imported ListOfPair from NMTDS;
    imported ListIteratorOfListOfPair  from NMTDS; 
 
    imported ListOfPairBoolean from NMTDS;
    imported ListIteratorOfListOfPairBoolean  from NMTDS; 
     
    imported ListOfIndexedDataMapOfShapeAncestorsSuccessors from NMTDS; 
    imported ListIteratorOfListOfIndexedDataMapOfShapeAncestorsSuccessors from NMTDS;  
    
    imported MapOfPassKey from NMTDS;
    imported MapIteratorOfMapOfPassKey from NMTDS; 
     
    imported MapOfPairBoolean from NMTDS;
    imported MapIteratorOfMapOfPairBoolean from NMTDS; 
    
    imported IndexedDataMapOfShapeBox from NMTDS;
    imported IndexedDataMapOfIntegerShape from NMTDS;
    imported IndexedDataMapOfShapeBndSphere from NMTDS;
 
    imported DataMapOfIntegerMapOfInteger from NMTDS;
    imported DataMapIteratorOfDataMapOfIntegerMapOfInteger from NMTDS;
     
    imported CArray1OfIndexRange from NMTDS;
	
end NMTDS;
