--  Copyright (C) 2007-2008  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
-- File:	NMTAlgo_Tools.cdl
-- Created:	Fri Jan 30 16:29:14 2004
-- Author:	Peter KURNEV
--		<pkv@irinox>


class Tools from NMTAlgo 

	---Purpose: 

uses  
    Orientation from TopAbs,

    Shape from TopoDS, 
    Edge  from TopoDS, 
    Face  from TopoDS,
    Shell from TopoDS, 
    	 
    ListOfShape from TopTools, 
    IndexedMapOfShape from TopTools
--raises

is
    OrientFacesOnShell (myclass; 
    	    aShell: Shell from TopoDS;  
	    aShellNew: out Shell from TopoDS); 
	 
    OrientFacesOnShell (myclass; 
    	    aF  : Face from TopoDS;  
	    aSh : out Shell from TopoDS);   
	    
    Orientation(myclass;  
    	    aE:  Edge from TopoDS; 
	    aF:  Face from TopoDS) 
	returns Orientation from TopAbs; 
	 
    Sense  (myclass;  
    	    aF1:  Face from TopoDS; 
	    aF2:  Face from TopoDS) 
	returns Integer from Standard; 
	 
    IsInside (myclass;  
    	    aS1:  Shape from TopoDS; 
    	    aS2:  Shape from TopoDS) 
    	returns Boolean from Standard;  
	 
    MakeShells(myclass; 
	aFC:Shape from TopoDS;
	aLS:out ListOfShape from TopTools);  
	
    MakeSolids(myclass; 
	aLS:out ListOfShape from TopTools);     

    MakeSolids(myclass; 
	aFC:Shape from TopoDS;
	aLS:out ListOfShape from TopTools);  
	 
    BreakWebs (myclass;  
    	    aS1:  Shape from TopoDS; 
    	    aS2:out Shape from TopoDS);  
	 
    FindImageSolid (myclass;  
    	    aFC  :  Shape from TopoDS;  
	    aMSo :  IndexedMapOfShape from TopTools;
    	    aSo  :  out Shape from TopoDS) 
    	returns Boolean from Standard;      
	    
--fields

end Tools;
