-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	NMTDS_Tools.cdl
--  Created:	Tue Feb 20 14:56:14 2007
--  Author:	Peter KURNEV
--
class Tools from NMTDS 

	---Purpose: 

uses
    ShapeEnum from TopAbs, 
    Vertex    from TopoDS,
    Shape     from TopoDS,
    IndexedDataMapOfShapeShape from TopTools 
    
--raises

is 
    TypeToInteger(myclass; 
    	    aT1: ShapeEnum from TopAbs; 
    	    aT2: ShapeEnum from TopAbs) 
    	returns Integer from Standard; 
	 
    HasBRep(myclass; 
    	    aT: ShapeEnum from TopAbs) 
    	returns Boolean from Standard;  
	 
    ComputeVV(myclass;  
    	    aV1:Vertex from TopoDS;  
    	    aV2:Vertex from TopoDS) 
    	returns Integer from Standard;  

    CopyShape(myclass; 
    	    aS:Shape from TopoDS;  
    	    aSC:out Shape from TopoDS);  

    CopyShape(myclass; 
    	    aS:Shape from TopoDS;  
    	    aSC  :out Shape from TopoDS; 
    	    aMSS :out IndexedDataMapOfShapeShape from TopTools);
--fields

end Tools;
