// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
//
-- File:	GEOMAlgo_PassKeyShape.cdl
-- Created:	
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 


class PassKeyShape from GEOMAlgo 
    inherits PassKey from GEOMAlgo  
    
	---Purpose: 

uses
    Shape from TopoDS, 
    ListOfShape from TopTools   
  	 
--raises

is 
    Create  
    	returns PassKeyShape from GEOMAlgo; 
      
    SetIds(me:out; 
    	    aS  :Shape from TopoDS); 
    	    
    SetIds(me:out; 
    	    aS1  :Shape from TopoDS; 
    	    aS2  :Shape from TopoDS); 
     
    SetIds(me:out; 
    	    aS1  :Shape from TopoDS; 
    	    aS2  :Shape from TopoDS; 
    	    aS3  :Shape from TopoDS); 
 
    SetIds(me:out;  
    	    aS1  :Shape from TopoDS; 
    	    aS2  :Shape from TopoDS; 
    	    aS3  :Shape from TopoDS;
    	    aS4  :Shape from TopoDS);
 
    SetIds(me:out;  
    	    aLS  :ListOfShape from TopTools); 
	     

fields 
    myUpper  : Integer from Standard is protected; 

end PassKeyShape;
