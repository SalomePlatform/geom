--  Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_BuilderTools.cdl
-- Created:	
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class BuilderTools from GEOMAlgo 

	---Purpose: 

uses
    Shape from TopoDS 

--raises

is 
    IsHole(myclass;  
    	    aW:  Shape from TopoDS;    
    	    aF:  Shape from TopoDS) 
	returns Boolean from Standard;

    IsHole(myclass;  
    	    aShell:  Shape from TopoDS)    
	returns Boolean from Standard;

--fields

end BuilderTools;
