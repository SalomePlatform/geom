--  Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_PassKey.cdl
-- Created:	Mon Nov 20 12:16:13 2006
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class PassKey from GEOMAlgo 

	---Purpose: 

uses
    Shape from TopoDS, 
    IndexedMapOfInteger from TColStd, 
    ListOfInteger from TColStd

--raises

is 
    Create  
    	returns PassKey from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_PassKey();" 
     
    Create(Other:PassKey from GEOMAlgo) 
    	returns PassKey from GEOMAlgo;
     
    Assign(me:out;  
    	    Other : PassKey from GEOMAlgo) 
    	returns PassKey from GEOMAlgo; 
    ---C++: alias operator =
    ---C++: return & 
	     
    Clear(me:out);
--    
    SetIds(me:out; 
    	    aI1  :Integer from Standard); 
	     
    SetIds(me:out; 
    	    aI1 :Integer from Standard; 
    	    aI2 :Integer from Standard);  
	     
    SetIds(me:out; 
    	    aI1 :Integer from Standard;    
    	    aI2 :Integer from Standard;    
    	    aI3 :Integer from Standard);  

    SetIds(me:out; 
    	    aI1 :Integer from Standard;    
    	    aI2 :Integer from Standard;    
    	    aI3 :Integer from Standard;    
    	    aI4 :Integer from Standard); 
     
    SetIds(me:out;  
    	    aLS  :ListOfInteger from TColStd);   

    NbIds(me) 
	returns Integer  from Standard; 
     
    IsEqual(me; 
    	    aOther:PassKey from GEOMAlgo) 
	returns Boolean from Standard;   		     
	 
    HashCode(me; 
	    Upper : Integer  from Standard)  
    	returns Integer from Standard;   	 
     
    Id(me; 
    	    aIndex: Integer  from Standard)  
    	returns  Integer from Standard;
    	

    Dump(me; 
    	aHex:Integer from Standard=0);  
     
	
fields 
    myNbIds: Integer from Standard is protected;  
    mySum  : Integer from Standard is protected;  
    myMap  : IndexedMapOfInteger from TColStd is protected; 

end PassKey;
