-- Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_Algo.cdl
-- Created:	Sat Dec 04 12:37:56 2004
-- Author:	Peter KURNEV
--		<peter@PREFEX>
--
deferred  class Algo from GEOMAlgo 

	---Purpose: 

--uses
--raises

is
    Initialize 
    	returns Algo from GEOMAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_Algo();" 

    Perform(me:out) 
	is deferred;      

    CheckData(me:out) 
	is virtual protected;  
    	
    CheckResult(me:out) 
	is virtual protected;
     
    ErrorStatus (me) 
    	returns Integer from Standard; 
  
    WarningStatus (me) 
    	returns Integer from Standard;

    ComputeInternalShapes(me : in out; theFlag : Boolean from Standard);
      ---Purpose: Allows to omit of creation of internal shapes (manifold topology).
      --          Needed for the SALOME/TRIPOLI module.

fields
    myErrorStatus   : Integer from Standard  is protected;	 
    myWarningStatus : Integer from Standard  is protected;	 
    myComputeInternalShapes : Boolean from Standard is protected;
 
end Algo;
