--  Copyright (C) 2007-2008  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
-- File:	NMTAlgo_Builder.cdl
-- Created:	Tue Jan 27 15:09:45 2004
-- Author:	Peter KURNEV
--		<pkv@irinox>


class Builder from NMTAlgo  
    inherits Algo from NMTAlgo 

	---Purpose: 

uses  
    Shape from TopoDS, 
    Face  from TopoDS,
    Edge  from TopoDS,
    IndexedMapOfShape                from TopTools, 
    IndexedDataMapOfShapeListOfShape from TopTools,  
    IndexedDataMapOfShapeShape       from TopTools,
    Image from BRepAlgo,
    DSFiller from NMTTools
--raises

is 
    Create 
    	returns Builder from NMTAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~NMTAlgo_Builder();" 

    Clear (me:out) 
    	is redefined;     	  
     
    ComputeWithFiller(me:out; 
    	aDSF: DSFiller from NMTTools) 
    	is redefined;  
     
    FillImagesEdges (me:out) 
    	is protected; 
	 
    FillIn2DParts (me:out) 
    	is protected; 
	 
    FillImagesFaces (me:out) 
    	is protected;  
	 
    FillSDFaces  (me:out) 
    	is protected; 
	
    ---  Queries 
    SplitVertices  (me:out) 
    	is protected;   

    IsSectionEdge (me;  
    	    E : Edge from TopoDS) 
        returns Boolean from Standard 
    	is protected;	  
	 
    HasSameDomainF(me;  
    	    F : Face from TopoDS)
        returns Boolean from Standard 
    	is protected;
    
    IsSameDomainF(me;  
    	    F1 : Face from TopoDS;
    	    F2 : Face from TopoDS)
        returns Boolean from Standard 
    	is protected;

fields 

    myImagesEdges       : Image from BRepAlgo is protected; 
    myImagesFaces       : Image from BRepAlgo is protected; 
    
    myQueryShapes       : IndexedMapOfShape                from TopTools is protected;
    -- 
    myIn2DParts         : IndexedDataMapOfShapeListOfShape from TopTools is protected;         
    mySectionParts      : IndexedDataMapOfShapeListOfShape from TopTools is protected; 
    mySDFaces           : IndexedDataMapOfShapeShape       from TopTools is protected;
    --	     
end Builder;
