// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
//
-- File:	GEOMAlgo_ShapeSolid.cdl
-- Created:	Thu Jan 13 12:44:07 2005
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2005


deferred class ShapeSolid from GEOMAlgo 
    	inherits Algo from GEOMAlgo 
	 
	---Purpose: 

uses 
    State from TopAbs,
    ListOfShape from TopTools, 
    PDSFiller from BOPTools,
    DSFiller  from BOPTools
--raises

is 
    Initialize 
    	returns ShapeSolid from GEOMAlgo;  
    

    SetFiller(me:out; 
    	    aDSF:DSFiller  from BOPTools); 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_ShapeSolid();"  
     
      
    Shapes(me;
	     aState:State from TopAbs) 
	returns ListOfShape from TopTools; 
    ---C++: return const &  
       
    BuildResult (me:out) 
	is deferred protected;	
    	
    Prepare(me:out)  
   	is deferred protected; 
	
fields
    myLSIN  :  ListOfShape from TopTools is protected;  
    myLSOUT :  ListOfShape from TopTools is protected;  
    myLSON  :  ListOfShape from TopTools is protected;  
    myRank  :  Integer from Standard is protected; 
    myDSFiller : PDSFiller from BOPTools is protected; 

end ShapeSolid;
