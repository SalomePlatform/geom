-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	NMTDS_Pair.cdl
--  Created:	
--  Author:	Peter KURNEV
--
class Pair from NMTDS 

	---Purpose: 

--uses
--raises

is 
    Create  
    	returns Pair from NMTDS; 
    ---C++: alias "Standard_EXPORT virtual ~NMTDS_Pair();" 

    Create(Other:Pair from NMTDS) 
    	returns Pair from NMTDS;
   ---C++: alias "Standard_EXPORT NMTDS_Pair& operator =(const NMTDS_Pair& Other);" 

    Clear(me:out);
	     
    SetIds(me:out; 
    	    aI1 :Integer from Standard; 
    	    aI2 :Integer from Standard);  
 
    Ids(me; 
    	    aI1 :out Integer from Standard;    
    	    aI2 :out Integer from Standard);	     
     
    IsEqual(me; 
    	    aOther:Pair from NMTDS) 
	returns Boolean from Standard;   		     
	 
    HashCode(me; 
	    Upper : Integer  from Standard)  
    	returns Integer from Standard;   	 
     
	
fields 
    myId1: Integer from Standard is protected;  
    myId2: Integer from Standard is protected;  

end Pair;
