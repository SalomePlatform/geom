--  Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
-- File:	GEOMAlgo_Tools.cdl
-- Created:	Mon Dec  6 11:26:02 2004
-- Author:	Peter KURNEV
--
class Tools from GEOMAlgo 

	---Purpose: 

uses    
    Pnt from gp, 
    Surface from Geom, 
    ShapeEnum from TopAbs,  
    Edge  from TopoDS, 
    Face  from TopoDS, 
    Shape from TopoDS,
    ListOfShape from TopTools,  
    IndexedDataMapOfShapeListOfShape from TopTools,
    Context from IntTools, 
    IndexedDataMapOfPassKeyShapeListOfShape from GEOMAlgo  --qft 
    
--raises

is   
    IsCompositeShape(myclass;  
    	    aS  :Shape from TopoDS) 
	returns Boolean from Standard;    

    RefineSDShapes(myclass; 
    	    aMSD:out IndexedDataMapOfPassKeyShapeListOfShape from GEOMAlgo; --qft
    	    aTol:Real from Standard; 
    	    aCtx:out Context from IntTools) 
    	returns Integer from Standard;

    FindSDShapes(myclass; 
    	    aLE :ListOfShape from TopTools;   
    	    aTol:Real from Standard; 
    	    aMEE:out IndexedDataMapOfShapeListOfShape from TopTools; 
	    aCtx:out Context from IntTools) 
    	returns Integer from Standard;
     
    FindSDShapes(myclass; 
    	    aE1   :Shape from TopoDS; 
	    aLE   :ListOfShape from TopTools; 
	    aTol  :Real from Standard;   
    	    aLESD :out ListOfShape from TopTools;
	    aCtx  :out Context from IntTools) 
    	returns Integer from Standard;  
	 
    ProjectPointOnShape(myclass;  
    	    aP1: Pnt from gp;  
    	    aS  :Shape from TopoDS;  
	    aP2:out Pnt from gp; 
    	    aCtx  :out Context from IntTools) 
        returns Boolean from Standard;  
  
    PointOnShape(myclass;  
    	    aS  :Shape from TopoDS; 
	    aP3D:out Pnt from gp); 
	     
    PointOnEdge(myclass;  
    	    aE  :Edge from TopoDS; 
	    aP3D:out Pnt from gp); 
	     
    PointOnEdge(myclass;  
    	    aE  :Edge from TopoDS; 
    	    aT  :Real from Standard;   
	    aP3D:out Pnt from gp); 

    PointOnFace(myclass;  
    	    aF  :Face from TopoDS; 
	    aP3D:out Pnt from gp); 
     
    PointOnFace(myclass;  
    	    aF  :Face from TopoDS; 
    	    aU  :Real from Standard; 
    	    aV  :Real from Standard; 
	    aP3D:out Pnt from gp);     

    RefinePCurveForEdgeOnFace  (myclass; 
    	    aE  :  Edge from TopoDS; 
            aF  :  Face from TopoDS; 
    	    aU1 : Real from Standard; 
    	    aU2 : Real from Standard); 

    IsUPeriodic(myclass;  
    	    aS:Surface from Geom) 
    	returns Boolean from Standard;   

    CorrectWires(myclass; 
    	    aS  :Shape from TopoDS) 
    	returns Boolean from Standard; 
--fields

end Tools;
