--  Copyright (C) 2007-2010  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_ClsfSolid.cdl
-- Created:	Mon Jan 29 10:28:07 2007
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class ClsfSolid from GEOMAlgo  
    inherits Clsf from GEOMAlgo 

	---Purpose: 

uses
    Shape from TopoDS
    
--raises

is
    Create 
    	returns mutable ClsfSolid from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_ClsfSolid();"  
      
    SetShape(me:mutable; 
    	    aS:Shape from TopoDS);  
	 
    Shape(me) 
    	returns Shape from TopoDS; 
    ---C++: return const &     
     
    Perform(me:mutable) 
	is redefined;      

    CheckData(me:mutable) 
	is redefined;  
    	 
    
fields  
    myShape: Shape from TopoDS is protected;
    myPClsf: Address from Standard is protected;
   
end ClsfSolid;
