--  Copyright (C) 2007-2008  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
--  File:	NMTDS_IndexRange.cdl
--  Created:	Fri Nov 28 10:31:05 2003
--  Author:	Peter KURNEV
--
class IndexRange from NMTDS 

	---Purpose: 

--uses
--raises

is 
    Create 
    	returns IndexRange from NMTDS; 
	 
    SetFirst(me:out; 
    	    aFirst:Integer from Standard);	 
	 
    SetLast(me:out; 
    	    aLast:Integer from Standard);	 
     
    First(me) 
    	returns Integer from Standard; 
	 
    Last(me) 
    	returns Integer from Standard; 				     

    IsInRange(me; 
    	    aIndex:Integer from Standard) 
    	returns Boolean from Standard; 

fields 
    myFirst  :  Integer from Standard is protected;  
    myLast   :  Integer from Standard is protected;  

end IndexRange;
