-- Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
-- 
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either 
-- version 2.1 of the License.
-- 
-- This library is distributed in the hope that it will be useful 
-- but WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public  
-- License along with this library; if not, write to the Free Software 
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
-- 
-- File:	NMTTools_PaveFiller.cdl
-- Created:	Fri Dec  5 14:35:00 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>


class PaveFiller from NMTTools 

	---Purpose: 

uses   
    DataMapOfIntegerInteger from TColStd,
    Pnt from gp,
    ShapeEnum  from  TopAbs, 
    Vertex     from  TopoDS, 
    Face       from  TopoDS,  
    Shape      from TopoDS, 
    -- Modified to add new definitions Thu Sep 14 14:35:18 2006 
    -- Contribution of Samtech www.samcef.com BEGIN 
    Edge       from  TopoDS, 
    ListOfShape from TopTools,  
    DataMapOfShapeShape from TopTools,
    ListOfInteger from TColStd,  
    -- Contribution of Samtech www.samcef.com END 
    
    Context     from IntTools, 
    ShrunkRange from IntTools,
    
    IndexedDataMapOfShapeInteger from BooleanOperations, 
    
    --InterferencePool  from BOPTools,
    --PInterferencePool from BOPTools, 
    PavePool          from BOPTools, 
    PaveBlock         from BOPTools,
    ListOfPaveBlock   from BOPTools,
    SplitShapesPool   from BOPTools, 
    Pave              from BOPTools, 
    PaveSet           from BOPTools, 
    Curve             from BOPTools, 
    SSInterference    from BOPTools, 
    
    IDMapOfPaveBlockIMapOfPaveBlock from BOPTools, 
    IDMapOfPaveBlockIMapOfInteger   from BOPTools, 
    SSIntersectionAttribute         from BOPTools, 
    
    CommonBlockPool         from NMTTools, 
    CommonBlock             from NMTTools, 
    ListOfCommonBlock       from NMTTools, 
   
    ShapesDataStructure  from NMTDS,  

    -- Modified to add new definitions Thu Sep 14 14:35:18 2006 
    -- Contribution of Samtech www.samcef.com BEGIN
    PShapesDataStructure from NMTDS, 
    Iterator             from NMTDS, 
    IndexedDataMapOfIndexedMapOfInteger from NMTTools,  
    -- Contribution of Samtech www.samcef.com END
     
    PIterator from NMTDS, 
    PInterfPool from NMTDS

--raises

is 
    Create 
    	returns PaveFiller from NMTTools;  
    ---C++: alias "Standard_EXPORT virtual ~NMTTools_PaveFiller();"
      
   -- Create(aIP:InterferencePool from BOPTools)
    --	returns PaveFiller from NMTTools; 
     
   -- Destroy (me: in out) 
	--is  virtual;    
    --  -C++: alias "Standard_EXPORT virtual ~NMTTools_PaveFiller(){Destroy();}"
    -- 
    --  Selectors/Modifiers
    --SetInterferencePool(me:out; 
    --	    aIP:PInterferencePool from BOPTools);
     
    SetCompositeShape (me:out;  
    	    aS:  Shape from TopoDS);  
     
    CompositeShape(me) 
    	returns  Shape from TopoDS; 
    	---C++:  return  const&  
	
    --InterfPool(me:out) 
    	--returns PInterferencePool from BOPTools; 

    --SetDS(me:out; 
    	--    aDS:PShapesDataStructure from NMTDS);  
	     
    DS(me:out) 
      	returns PShapesDataStructure from NMTDS;  
     
    --SetDSIt(me:out; 
    	--    	aIt:PIterator from NMTDS); 
	 
    DSIt(me:out) 
    	returns PIterator from NMTDS; 
     
    IP(me:out)  
    	returns PInterfPool from NMTDS; 
    --	 
    --  Perform the algo  
    -- Modified to add new method Thu Sep 14 14:35:18 2006 
    -- Contribution of Samtech www.samcef.com BEGIN      
    Init       (me:out) 
    	is virtual  protected; 
    -- Contribution of Samtech www.samcef.com END
	 
    Clear   (me:out) 
    	is virtual  protected;

    Perform    (me:out) 
	is virtual;   
	 
    PerformVV  (me:out) 
    	is virtual protected;  
     
    PerformVE  (me:out) 
    	is virtual protected; 
     
    PerformVF  (me:out) 
    	is virtual protected; 

    PerformEE (me:out) 
    	is virtual protected; 
      
    PerformEF (me:out) 
    	is virtual protected; 
   
    PerformFF (me:out) 
    	is virtual protected; 
     
    MakeSplitEdges(me:out) 
    	is protected;   
     
    PreparePaveBlocks (me:out; 
    	    aType1: ShapeEnum  from  TopAbs; 
    	    aType2: ShapeEnum  from  TopAbs) 
    	is virtual protected; 
     
    CorrectShrunkRanges(me:out; 
    	    aSide:  Integer  from  Standard; 
    	    aPave:  Pave from BOPTools; 
    	    aSR  :  out ShrunkRange  from  IntTools)
    	is protected; 
	 
    PreparePaveBlocks (me:out;   
    	    anE:Integer from Standard) 
    	is virtual protected;  		  
		       
    --PerformNewVertices  (me:out) 
    	--is virtual;  
     
    PrepareEdges  (me:out) 
    	is virtual protected;  
     
    --SortTypes      (me;   
    --	    anInd1:in out Integer from Standard; 
    --        anInd2:in out Integer from Standard) 
    --	is protected; 
     
    --ExpectedPoolLength(me) 
    --	returns  Integer from Standard 
	--is protected;  
    --
    -- Query section 
    IsDone(me) 
    	returns  Boolean from Standard; 

    Context(me) 
    	 returns Context from IntTools; 
    	---C++:return const &	

    ChangeContext(me:out) 
    	 returns Context from IntTools;  
    	---C++:return &	

    PavePool(me) 
    	returns  PavePool from BOPTools; 
    	---C++:return const &	 

    ChangePavePool(me:out) 
    	returns  PavePool from BOPTools; 
    	---C++:return &	

    CommonBlockPool(me) 
    	returns  CommonBlockPool from NMTTools; 
    	---C++:return const &	 

    ChangeCommonBlockPool(me:out) 
    	returns  CommonBlockPool from NMTTools; 
    	---C++:return &	

    SplitShapesPool(me)  
    	returns  SplitShapesPool from BOPTools;
    	---C++:return const &	

    ChangeSplitShapesPool(me:out)  
    	returns  SplitShapesPool from BOPTools;
    	---C++:return  &	
     
    FindSDVertex (me; 
    	    	    nV:  Integer  from  Standard) 
    	returns Integer from Standard; 

    IsSuccessorsComputed (me;  
    	    iF1:Integer from  Standard; 
    	    iF2:Integer from  Standard) 
    	returns  Boolean from Standard 
    	is protected;  

    IsBlocksCoinside (me; 
    	    aPB1:PaveBlock from BOPTools;
    	    aPB2:PaveBlock from BOPTools) 
	returns Boolean from Standard 
    	is protected; 
     
    RefinePavePool(me:out) 
    	is protected;  

    CheckFacePaves(me:out;  
    	     aV : Vertex  from TopoDS;  
     	     nF:  Integer from Standard) 
    	returns Integer from Standard 
    	is protected;  
	 
    ReplaceCommonBlocks (me:out; 
	    aLCB: ListOfCommonBlock from NMTTools) 
        is protected; 
     
    RemoveCommonBlocks (me:out; 
	    aLCB: ListOfCommonBlock from NMTTools) 
        is protected;
     
    SplitCommonBlocks (me:out; 
	    aLCB: ListOfCommonBlock from NMTTools) 
        is protected;  

    SplitCommonBlock (me:out; 
    	    aCB : CommonBlock from NMTTools; 
	    aLCB: out ListOfCommonBlock from NMTTools) 
        is protected; 

    EECommonBlocks(me:out; 
    	    aM:IDMapOfPaveBlockIMapOfPaveBlock from BOPTools) 
    	is protected; 
     
    EFCommonBlocks(me:out;  
    	     aMapCB:IDMapOfPaveBlockIMapOfInteger from BOPTools) 
        is protected;  
	 
    EENewVertices (me:out;  
    	    aM:IndexedDataMapOfShapeInteger from BooleanOperations) 
    	is protected;  

    EENewVertices (me:out;  
    	    aV:Vertex from TopoDS;  
    	    aM:IndexedDataMapOfShapeInteger from BooleanOperations) 
    	is protected; 
     
    EFNewVertices (me:out; 
    	    aM:IndexedDataMapOfShapeInteger from BooleanOperations) 
    	is protected; 
     
    EFNewVertices (me:out; 
    	    aV:Vertex from TopoDS;  
    	    aM:IndexedDataMapOfShapeInteger from BooleanOperations) 
    	is protected;   
	 
    UpdateCommonBlocks(me:out) 
    	is protected;  
     
    UpdatePaveBlocks(me:out) 
    	is protected; 
	 
    SplitIndex(me; 
    	    aPB:PaveBlock from BOPTools) 
	returns Integer from Standard  
    	is protected;		     
    	 
    MakeBlocks(me:out) 
    	is protected;   

    -------------------------------------------------------------- 
    ---	  
    ---  Some API FUNCTIONS  
    ---  	    	 
    SplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  

    SplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	
    SplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	
    SplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	
    SplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	
    SplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
     
    SplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
     
    SplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
     
    SplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  

    SplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
    --
    SplitsFace  (me:out;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  

    SplitsFace  (me:out;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  

    CommonBlocksFace (me:out;  
    	         nF  :Integer from Standard;  
    	         aLCB:out ListOfCommonBlock from NMTTools) 
    	returns Integer from Standard;   
	
    PrepareFace(me:out;  
    	    nF  :  Integer from Standard; 
    	    aF  : out Face from TopoDS); 
     
    -- 
    RealPaveBlock(me:out;   
    	    aPB:PaveBlock from BOPTools) 
	returns PaveBlock from BOPTools; 
    ---C++: return const & 	  
    
    -- Modified to add new method Thu Sep 14 14:35:18 2006 
    -- Contribution of Samtech www.samcef.com BEGIN  
    RealPaveBlock(me:out;   
    	    aPB:PaveBlock from BOPTools; 
    	    aLB:out ListOfInteger from TColStd) 
	returns PaveBlock from BOPTools; 
    ---C++: return const & 	 
    -- Contribution of Samtech www.samcef.com END 
     
    RealSplitsFace  (me:out;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
	 
    HasRealSplitsInOnFace (me:out; 
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard) 
    	returns Boolean from Standard; 
	 
    RealSplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
     
    RealSplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
     
    RealSplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
     
    RealSplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 

    RealSplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
    --   
    PrepareSetForFace(me:out;   
    	    	nF1 :Integer from Standard;  
    	        nF2 :Integer from Standard;  
		aLPB: ListOfPaveBlock from BOPTools;  
    	    	aPSF:out PaveSet from BOPTools); 
		 
    PutPaveOnCurve(me:out;   
    	    	aPSF: PaveSet from BOPTools; 
		aTol: Real from Standard;  
		aBC : out Curve from BOPTools); 
	 
    PutBoundPaveOnCurve (me:out; 
    	    	    aBC :out Curve from BOPTools;	 
     	    	    aFF :out SSInterference from BOPTools); 
    	
    PutBoundPaveOnCurve (me:out;  
    	    	    aP  : Pnt from  gp; 
		    aT  : Real from Standard; 			 
    	    	    aBC :out Curve from BOPTools;	 
     	    	    aFF :out SSInterference from BOPTools); 
    	
    FindPave            (me:out; 
		    aP  : Pnt from gp;  
    	    	    aTpV: Real from Standard;  
    	    	    aPS : PaveSet from BOPTools; 
		    aPV :out Pave from BOPTools) 
    	returns Boolean from Standard; 
	 
    CheckIntermediatePoint(me:out;  
    	    	    aPB : PaveBlock      from BOPTools;  
    	    	    aPBR: PaveBlock      from BOPTools;  
     	    	    aTol: Real  from  Standard) 
    	returns Integer from Standard; 	
		

    IsExistingPaveBlock (me:out; 
    	    	    aPB : PaveBlock       from BOPTools; 
     	    	    aLPB: ListOfPaveBlock from BOPTools; 
    	    	    aTol: Real  from  Standard) 
    	returns Boolean from Standard;  
	  
    MakePCurves (me:out); 
     
    -- Modified to add new methods Thu Sep 14 14:35:18 2006 
    -- Contribution of Samtech www.samcef.com BEGIN
    PerformVF1(me:out) 
    	is protected;  
	 
    MakeAloneVertices(me:out) 
    	is protected;   
	 
    AloneVertices(me)  
    	returns IndexedDataMapOfIndexedMapOfInteger from NMTTools; 
    ---C++: return const & 
    -- Contribution of Samtech www.samcef.com END 
     
    IsExistingPaveBlock (me:out; 
    	    	    aPB : PaveBlock   from BOPTools; 
     	    	    aLPB: ListOfShape from TopTools; 
    	    	    aTol: Real  from  Standard) 
    	returns Boolean from Standard;  

    --
    CheckCoincidence (me:out; 
    	    	    aPB : PaveBlock   from BOPTools; 
     	    	    aLPB: ListOfPaveBlock from BOPTools) 
    	returns Boolean from Standard;  
    -- 
     
    CheckIntermediatePoint(me:out;  
    	    	    aPB : PaveBlock      from BOPTools;  
    	    	    aE  : Edge from TopoDS;  
     	    	    aTol: Real  from  Standard) 
    	returns Integer from Standard; 	 

    -- Modified to add new method Thu Sep 14 14:35:18 2006 
    -- Contribution of Samtech www.samcef.com BEGIN
    SharedEdges(me:out;  
    	         nF1  :Integer from Standard;  
    	         nF2  :Integer from Standard;  
    	         aLNE :out ListOfInteger from TColStd; 
    	         aLSE :out ListOfShape   from TopTools); 
    -- Contribution of Samtech www.samcef.com END 

    FuseVertices(me; 
    	aC:Shape from TopoDS; 
	aDMVV:  out  DataMapOfShapeShape from TopTools);  
     
fields 
    --myIntrPool         :  PInterferencePool from BOPTools    	is protected; 
    myDS               :  PShapesDataStructure from NMTDS   	is protected;   
    myIsDone           :  Boolean from Standard                 is protected; 
    myNbSources        :  Integer from Standard                 is protected;  
    myNbEdges          :  Integer from Standard           	is protected;  

    myPavePool         :  PavePool from BOPTools                is protected;     
    myPavePoolNew      :  PavePool from BOPTools                is protected;  
    myCommonBlockPool  :  CommonBlockPool from NMTTools         is protected;  
    mySplitShapesPool  :  SplitShapesPool from BOPTools	        is protected;    
    -- 
    myContext          :  Context from IntTools                 is protected; 
    mySectionAttribute :  SSIntersectionAttribute from BOPTools is protected; 
    myAloneVertices    :  IndexedDataMapOfIndexedMapOfInteger from NMTTools is protected;   
    --modified by NIZNHY-PKV Wed Oct 11 11:06:50 2006f
    myVSD              :  DataMapOfIntegerInteger from TColStd is protected; 
    myDSIt             :  PIterator from NMTDS is protected;  
    myCompositeShape   :  Shape from TopoDS is protected;
    myIP               :  PInterfPool from NMTDS is protected;     
    --modified by NIZNHY-PKV Wed Oct 11 11:06:55 2006t 
end PaveFiller;
