-- File:	NMTTools_DEProcessor.cdl
-- Created:	Wed Sep 12 12:08:37 2001
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2001


class DEProcessor from NMTTools 

	---Purpose:  
    	--   
    	--  The  Algorithm to compute and store in interferences' pool 
	--- and in the Data  Structure  the following values        
    	--- for degenerated edges 
	---         1.  Paves/Pave set(s)
	---         2.  Split parts 
	---         3.  States (3D) for split parts 
        --- 
	
uses  

    Vertex from TopoDS,
    Edge   from TopoDS, 
    Face   from TopoDS, 
     
    PPaveFiller     from NMTTools, 
    PaveFiller      from NMTTools, 
    --PDSFiller       from NMTTools,   
    ListOfPaveBlock from BOPTools,
    PShapesDataStructure from NMTDS, 
    IndexedDataMapOfIntegerDEInfo from BOPTools	  


is
    --Create (aFiller:out PDSFiller from NMTTools) 
    --	returns  DEProcessor from NMTTools; 
    	---Purpose:  
    	--- Constructor 
    	--- 
    Create (aFiller:out PaveFiller from NMTTools) 
    	returns  DEProcessor from NMTTools; 
    	---Purpose:  
    	--- Constructor 
    	---	
    Do(me:out);   
    	---Purpose: 
    	--- Launches the processor   
    	---
    IsDone(me) 
    	returns Boolean from Standard; 
    	---Purpose:  
    	--- Returns TRUE if it is Ok       
    	---
    --- 
    ---    Private block 
    ---
    ---
    FindDegeneratedEdges (me:out) 
    	is  protected; 
	
    DoPaves  (me:out) 
    	is  protected; 
	 
    FindPaveBlocks (me:out; 
    	    nED:Integer from Standard; 
    	    nVD:Integer from Standard; 
    	    nFD:Integer from Standard; 
    	    aLPB:out ListOfPaveBlock from BOPTools) 
    	is  protected; 
     
    FillPaveSet (me:out; 
    	    nED:Integer from Standard; 
    	    nVD:Integer from Standard; 
    	    nFD:Integer from Standard; 
    	    aLPB: ListOfPaveBlock from BOPTools) 
    	is  protected; 

    FillSplitEdgesPool(me:out; 
    	    nED:Integer from Standard)
    	is  protected; 
  
    MakeSplitEdges(me:out; 
    	    nED:Integer from Standard;
    	    nFD:Integer from Standard)
    	is  protected;   
	 
    MakeSplitEdge  (me:out;   
        	    aS1: Edge from TopoDS; 
		    aF : Face from TopoDS;	     
		    aV1: Vertex from TopoDS;	     
   	    	    aP1: Real from Standard; 
    	    	    aV2: Vertex from TopoDS; 
		    aP2: Real from Standard; 
    	    	    aNewEdge:out Edge from TopoDS) 
    	is protected; 		
     
fields 
        
    --myDSFiller: PDSFiller   from NMTTools is protected;
    myFiller  : PPaveFiller from NMTTools is protected; 
    myDS      : PShapesDataStructure from NMTDS is protected;
    myIsDone  : Boolean   from Standard is protected;   
    myDEMap   : IndexedDataMapOfIntegerDEInfo from BOPTools is protected; 
	     
end DEProcessor;
