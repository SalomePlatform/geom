--  Copyright (C) 2007-2010  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_BuilderSolid.cdl
-- Created:	
-- Author:	Peter KURNEV  
--
class BuilderSolid from GEOMAlgo 
    	inherits BuilderArea from GEOMAlgo 
	 
	---Purpose: The algorithm to build solids from set of faces  

--uses 
--raises

is 
    Create  
    	---Purpose:  Empty  constructor
    	returns BuilderSolid from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_BuilderSolid();" 
     
     
    Perform(me:out)  
    	---Purpose:  Performs the algorithm 
    	is redefined;  
	 
    PerformShapesToAvoid(me:out) 
	---Purpose:  Collect the faces that 
	--           a) are internal        	 
	--           b) are the same and have different orientation         	 
    	is redefined protected; 
	 
    PerformLoops(me:out) 
	---Purpose: Build draft shells 
        --          a)myLoops - draft shells that consist of  
        --                       boundary faces 
	--          b)myLoopsInternal - draft shells that contains 
	--                               inner faces 
    	is redefined protected;  
	 
    PerformAreas(me:out)   
    	---Purpose: Build draft solids that contains boundary faces   
    	is redefined protected;  

    PerformInternalShapes(me:out)   
    	---Purpose: Build finalized solids with internal shells   
    	is redefined protected;   

--fields 
  
end BuilderSolid; 
