// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
// See http://www.salome-platform.org/
//
--  GEOM PARTITION : partition algorithm
--
--  Copyright (C) 2003  CEA/DEN, EDF R&D
--
--
--
--  File   : Partition_Loop2d.cdl
--  Author : Benedicte MARTIN
--  Module : GEOM

class Loop2d from Partition

        ---Purpose: Builds the loops from a set of edges on a face.
	--          It works in  supposition  that  all constant edges
	--          are split edges of  an initialization face and all
	--          section edges are new on the face

uses

    Orientation               from TopAbs,
    Boolean                   from Standard,
    Face                      from TopoDS,
    Image                     from BRepAlgo,
    Face                      from TopoDS,
    Edge                      from TopoDS,
    ListOfShape               from TopTools,
    DataMapOfShapeListOfShape from TopTools,
    MapOfShape                from TopTools
is

    Create;
    
    Init (me : in out; F : Face from TopoDS)
	---Purpose: Init with <F> the set of edges must have
	--          pcurves on <F>. 
    is static;
    
    AddConstEdge  (me : in out; E : Edge from TopoDS)
	---Purpose: Add <E> as unique edge in the result.
    is static;

    AddSectionEdge  (me : in out; E : Edge from TopoDS)
	---Purpose: Add <E> as double edge in the result.
    is static;

    Perform(me : in out)
	---Purpose: Make loops.
    is static;
    
    NewWires (me)	
	---Purpose: Returns the list of wires performed. 
	--          can be an empty list.
	---C++: return const &
    returns ListOfShape from TopTools;
    	
    WiresToFaces (me : in out; EdgeImage : Image      from BRepAlgo)
    	---Purpose:  Build faces from the wires result.
    	--           <EdgeImage> serves to  find  original edge by new
    	--           one.
    is static;
    
    NewFaces (me)
        ---Purpose: Returns the list of faces.
    	---Warning: The method <WiresToFaces> as to be called before.
    	--          can be an empty list.
	---C++: return const &
    returns ListOfShape from TopTools;

    
fields

    myFace       : Face        from TopoDS;
    myFaceOri    : Orientation from TopAbs;
    myConstEdges : ListOfShape from TopTools;
    myNewWires   : ListOfShape from TopTools;
    myNewFaces   : ListOfShape from TopTools;

     -- internal wires do not contain constant edges
    myInternalWL : ListOfShape from TopTools;
    
    mySectionEdges : MapOfShape from TopTools;
    
end Loop2d;
