-- Copyright (C) 2006 SAMTECH 
-- 
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either 
-- version 2.1 of the License.
-- 
-- This library is distributed in the hope that it will be useful 
-- but WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public  
-- License along with this library; if not, write to the Free Software 
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
-- 
-- File:	NMTDS_PassKeyBoolean.cdl
-- Created:	
-- Author:	Peter KURNEV
--		<pkv@irinox>


class PassKeyBoolean from NMTDS 
    inherits  PassKey from NMTDS 

	---Purpose: 

uses
    Shape from TopoDS, 
    ListOfInteger from TColStd   
  	 
--raises

is 
    Create  
    	returns PassKeyBoolean from NMTDS; 
     
    Assign(me:out;  
    	    Other : PassKeyBoolean from NMTDS) 
    	returns PassKeyBoolean from NMTDS; 
    ---C++: alias operator =
    ---C++: return & 
--     
    SetFlag(me:out; 
    	    aFlag: Boolean from Standard); 
	 
    Flag(me)  
    	returns Boolean from Standard;      

fields 
 
    myFlag: Boolean from Standard is protected;  

end PassKeyBoolean;
