--  Copyright (C) 2007-2010  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	BlockFix_SphereSpaceModifier.cdl
--  Created:	Tue Dec  7 12:01:49 2004
--  Author:	Pavel Durandin
--
class SphereSpaceModifier from BlockFix inherits Modification from BRepTools 

	---Purpose: Rotation of the parametric space of the sphere in order
        --          to avoid the seam and degenerared edge within it

uses
    Vertex   from TopoDS, 
    Edge     from TopoDS,
    Face     from TopoDS,
    Location from TopLoc,
    Shape    from GeomAbs,
    Pnt      from gp,
    Curve    from Geom,
    Curve    from Geom2d,
    Surface  from Geom,
    IndexedMapOfTransient from TColStd,
    DataMapOfShapeInteger from TopTools

is
    
    Create returns mutable SphereSpaceModifier from BlockFix;
    
    SetTolerance(me: mutable; Toler: Real);
    	---Purpose: Sets the tolerance for recognition of geometry

    NewSurface(me: mutable; F  :     Face     from TopoDS;
                            S  : out Surface  from Geom;
		            L  : out Location from TopLoc;
		            Tol: out Real     from Standard;
                            RevWires : out Boolean from Standard;
                            RevFace  : out Boolean from Standard)
    returns Boolean from Standard;
      	---Purpose: Returns Standard_True if the face <F> has  been
	--          modified. In this case, <S> is the new geometric
	--          support of the face, <L> the new location,  <Tol>
	--          the new tolerance.  Otherwise, returns
	--          Standard_False, and <S>, <L>, <Tol> are  not
	--          significant.
	
    NewCurve(me: mutable; E  :     Edge     from TopoDS;
                          C  : out Curve    from Geom;
		          L  : out Location from TopLoc;
		          Tol: out Real     from Standard)
    returns Boolean from Standard;
	---Purpose: Returns Standard_True  if  the edge  <E> has  been
	--          modified.  In this case,  <C> is the new geometric
	--          support of the  edge, <L> the  new location, <Tol>
	--          the         new    tolerance.   Otherwise, returns
	--          Standard_False,    and  <C>,  <L>,   <Tol> are not
	--          significant.

    NewPoint(me: mutable; V  :     Vertex   from TopoDS;
                          P  : out Pnt      from gp;
		          Tol: out Real     from Standard)
    returns Boolean from Standard;
	---Purpose: Returns  Standard_True if the  vertex <V> has been
	--          modified.  In this  case, <P> is the new geometric
	--          support of the vertex,   <Tol> the new  tolerance.
	--          Otherwise, returns Standard_False, and <P>,  <Tol>
	--          are not significant.

    NewCurve2d(me: mutable; E    :     Edge     from TopoDS;
                            F    :     Face     from TopoDS;
                            NewE :     Edge     from TopoDS;
                            NewF :     Face     from TopoDS;
                            C    : out Curve    from Geom2d;
		            Tol  : out Real     from Standard)
    returns Boolean from Standard;
    	---Purpose: Returns Standard_True if  the edge  <E> has a  new
	--          curve on surface on the face <F>.In this case, <C>
	--          is the new geometric support of  the edge, <L> the
	--          new location, <Tol> the new tolerance.
	--          
	--          Otherwise, returns  Standard_False, and <C>,  <L>,
	--          <Tol> are not significant.
	--          
	--          <NewE> is the new  edge created from  <E>.  <NewF>
	--          is the new face created from <F>. They may be usefull.

    NewParameter(me: mutable; V  :     Vertex from TopoDS;
                              E  :     Edge   from TopoDS;
                              P  : out Real   from Standard;
  		              Tol: out Real   from Standard)
    returns Boolean from Standard;
	---Purpose: Returns Standard_True if the Vertex  <V> has a new
	--          parameter on the  edge <E>. In  this case,  <P> is
	--          the parameter,    <Tol>  the     new    tolerance.
	--          Otherwise, returns Standard_False, and <P>,  <Tol>
	--          are not significant.

    Continuity(me: mutable; E          : Edge from TopoDS;
    	                    F1,F2      : Face from TopoDS;
			    NewE       : Edge from TopoDS;
			    NewF1,NewF2: Face from TopoDS)
    returns Shape from GeomAbs;
	---Purpose: Returns the  continuity of  <NewE> between <NewF1>
	--          and <NewF2>.
	--          
	--          <NewE> is the new  edge created from <E>.  <NewF1>
	--          (resp. <NewF2>) is the new  face created from <F1>
	--          (resp. <F2>).
    
    ForRotation(me: mutable; F: Face from TopoDS) returns Boolean;
    
fields 
    
    myTolerance   : Real;
    myMapOfFaces  : DataMapOfShapeInteger from TopTools;
    myMapOfSpheres: IndexedMapOfTransient from TColStd;
    --myMapOfGeom: MapOfShapeTransient from TColStd;

end SphereSpaceModifier;

