-- File:	BlockFix_BlockFixAPI.cdl
-- Created:	Tue Dec  7 17:56:09 2004
-- Author:	Pavel Durandin
--		<det@doomox>
---Copyright:	Open CASCADE SA 2004

class BlockFixAPI from BlockFix inherits TShared from MMgt

	---Purpose: 

uses

    Shape from TopoDS,
    ReShape from ShapeBuild 

is
    Create returns BlockFixAPI from BlockFix;
    	---Purpose: Empty constructor
	
    SetShape(me: mutable; Shape: Shape from TopoDS);
    	---Purpose: Sets the shape to be operated on
	---C++: inline

    Perform(me: mutable);
    	---Purpose: 
	
    Shape(me) returns Shape from TopoDS;
    	---Purpose: Returns resulting shape.
	---C++: inline
    
    Context(me:mutable) returns ReShape from ShapeBuild;
    	---Purpose: Returns modifiable context for storing the 
	--          mofifications
	---C++: inline
    	---C++: return &
    
    Tolerance (me:mutable) returns Real;
    	---Purpose: Returns modifiable tolerance of recognition
    	---C++: inline
    	---C++: return &

fields
    
    myContext     : ReShape from ShapeBuild;
    myShape       : Shape from TopoDS;
    myTolerance   : Real from Standard;
  
end BlockFixAPI from BlockFix;
