--  GEOM GEOMDS : implementation of Geometry component data structure and Geometry documents management
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : GEOMDS_Application.cdl
--  Author : Yves FRICAUD
--  Module : GEOM

class Application from GEOMDS  inherits Application from TDocStd

	---Purpose: 

uses
    Label                    from TDF,
    SequenceOfExtendedString from TColStd,
    CString                  from Standard,
    Document                 from TDocStd


is

    Create 
    returns mutable Application from GEOMDS;
    
    Formats(me: mutable; Formats: out SequenceOfExtendedString from TColStd) 
    is redefined;    

    ResourcesName (me: mutable) returns CString from Standard;

end Application;
