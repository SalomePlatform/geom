// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
// See http://www.salome-platform.org/
//
-- File:	GEOMAlgo_FinderShapeOn1.cdl
-- Created:	Fri Mar  4 10:26:54 2005
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2005


class FinderShapeOn1 from GEOMAlgo  
    inherits ShapeAlgo from GEOMAlgo 

	---Purpose: 

uses
    Surface from Geom, 
    Surface from GeomAdaptor, 
     
    ShapeEnum from TopAbs, 
    State from TopAbs,
    Face from TopoDS, 
    Edge from TopoDS, 
    ListOfShape from TopTools,  
     
    State from GEOMAlgo, 
    ListOfPnt from GEOMAlgo, 
    IndexedDataMapOfShapeState from GEOMAlgo 
    
--raises

is 
    Create   
    	returns FinderShapeOn1 from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_FinderShapeOn1();" 

    SetSurface(me:out; 
    	    aS:Surface from Geom); 
	 
    SetShapeType(me:out; 
    	    aST:ShapeEnum from TopAbs); 
	 
    SetState(me:out; 
    	    aSF:State from GEOMAlgo);      
     
    SetNbPntsMin(me:out; 
    	    aNb:Integer from Standard);   

    NbPntsMin(me) 
    	returns Integer from Standard; 
	 
    SetNbPntsMax(me:out; 
    	    aNb:Integer from Standard);   

    NbPntsMax(me) 
    	returns Integer from Standard; 
	 
    Surface(me) 
    	returns Surface from Geom; 
    ---C++: return const & 
     
    ShapeType(me) 
    	returns ShapeEnum from TopAbs; 
	 
    State(me)
    	returns State from GEOMAlgo;  
     
    Perform(me:out) 
	is redefined; 
    	 
    Shapes(me)
	returns ListOfShape from TopTools; 
    ---C++: return const &  
    -- 
    --  protected  methods
    -- 
    CheckData(me:out) 
	is redefined protected; 
	 
    ProcessVertices(me:out) 
    	is protected; 
     
    ProcessEdges(me:out) 
    	is protected; 
  
    ProcessFaces(me:out) 
    	is protected; 
	 
    ProcessSolids(me:out) 
    	is protected; 
	  
    InnerPoints(me:out; 
	    aF :Face from TopoDS;   	     
    	    aLP:out ListOfPnt from GEOMAlgo) 
    	is protected;  
	 
    InnerPoints(me:out; 
	    aE :Edge from TopoDS;   	     
    	    aLP:out ListOfPnt from GEOMAlgo) 
    	is protected; 
	 
    InnerPoints(me:out; 
	    aE :Edge from TopoDS;   	     
	    aNbPnts: Integer from Standard;     
	    aLP:out ListOfPnt from GEOMAlgo) 
    	is protected;  
      
    MSS (me)  
    	returns IndexedDataMapOfShapeState from GEOMAlgo; 
    ---C++:return const &  	
    
    GetPointState(me:out; aP: Pnt from gp)
        returns State from TopAbs is virtual protected;

fields
    mySurface   : Surface from Geom is protected;  
    myShapeType : ShapeEnum from TopAbs is protected;  
    myState     : State from GEOMAlgo is protected;  
    myNbPntsMin : Integer from Standard is protected;   
    myNbPntsMax : Integer from Standard is protected;   
    -- 
    myGAS       : Surface from GeomAdaptor is protected;
    myLS        : ListOfShape from TopTools is protected; 
    --     
    myMSS       : IndexedDataMapOfShapeState from GEOMAlgo is protected;
 
end FinderShapeOn1;
