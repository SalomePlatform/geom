-- File:	Partition_Loop3d.cdl
-- Created:	Mon Oct 21 09:47:19 2002
---Copyright:	 OPEN CASCADE 2002

class Loop3d from Partition

        ---Purpose: Builds the shells from a set of faces.
        --          Provides  methods   for   comparing  faces  mutual
        --          location.
        
uses
    Vec                              from gp,
    MapOfOrientedShape               from TopTools,
    IndexedDataMapOfShapeListOfShape from TopTools,
    Face                             from TopoDS,
    Edge                             from TopoDS,
    ListOfShape                      from TopTools,
    Shape                            from TopoDS
    
is

    Create;
    
    AddConstFaces  (me : in out; S : Shape from TopoDS)
	---Purpose: Add faces of <S> as unique faces in the result.
    is static;

    AddSectionFaces  (me : in out; S : Shape from TopoDS)
	---Purpose: Add faces of <S> as double faces in the result.
    is static;

    MakeShells (me : in out; AvoidFacesMap : MapOfOrientedShape from TopTools)
        returns ListOfShape from TopTools is static;
        ---Purpose: Make and return shells. 
        --          <AvoidFacesMap> can contain faces that must not be
        --          added to result shells.
        ---C++: return const &
    
    
        ---Category: class methods
    
    IsInside (myclass; E        : Edge    from TopoDS;
                       F1, F2   : Face    from TopoDS;
                       CountDot : Boolean from Standard;
                       Dot      : in out Real    from Standard;
                       GoodOri  : in out Boolean from Standard)
        returns Boolean from Standard;
        ---Purpose: check if <F2> is inside <F1> by edge <E>.
        --          if <CountDot>, compute <Dot>: scalar production of
        --          normalized  vectors  pointing  inside  faces,  and
        --          check if faces are oriented well for sewing
    
    Normal (myclass; E : Edge from TopoDS;
                     F : Face from TopoDS) returns Vec from gp;
    
    
fields

    myNewShells : ListOfShape from TopTools; -- result
    
    myFaces     : ListOfShape from TopTools;
    myEFMap     : IndexedDataMapOfShapeListOfShape from TopTools;
    
end Loop3d;
