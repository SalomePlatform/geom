-- File:	GEOMAlgo.cdl
-- Created:	Sat Dec 04 12:36:22 2004
-- Author:	Peter KURNEV
--		<peter@PREFEX>
---Copyright:	 Matra Datavision 2004


package GEOMAlgo 

	---Purpose: 

uses  
    TCollection, 
    TColStd, 
    Geom,     
    Bnd, 
    gp,	 
    TopAbs,
    TopoDS, 
    TopTools, 
    IntTools, 
    BOPTools, 
    BOP     
    
is   
    --  enumerations 
    --
    enumeration State is 
    	ST_UNKNOWN, 
	ST_IN,
	ST_OUT,
	ST_ON, 
	ST_ONIN, 
	ST_ONOUT, 
	ST_INOUT    
    end State;
    -- 
    --  classes 
    -- 
    deferred class Algo;
    deferred class ShapeAlgo; 
    -- 
    --  gluer    	     
    class Gluer; 
    class GlueAnalyser; 
    class CoupleOfShapes; 
    class PassKey; 
    class PassKeyMapHasher; 
    class SurfaceTools; 
    class Tools; 
    --	     
    --  finder on 
    deferred class ShapeSolid;
    class WireSolid; 
    class ShellSolid; 
    class VertexSolid; 
    class SolidSolid; 
    class FinderShapeOn; 
    --
    --  instantiations
    class IndexedDataMapOfPassKeyListOfShape   
	instantiates IndexedDataMap from TCollection (PassKey from GEOMAlgo, 
						      ListOfShape from TopTools, 
                                                      PassKeyMapHasher from GEOMAlgo); 
     
    class IndexedDataMapOfShapeBox  
    	instantiates IndexedDataMap from TCollection   	(Shape from TopoDS,
	    		    		         	 Box from Bnd,
	    		    		         	 ShapeMapHasher from TopTools);
    class IndexedDataMapOfIntegerShape  
    	instantiates IndexedDataMap from TCollection   	(Integer from Standard,
	    		    		         	 Shape from TopoDS,
	    		    		         	 MapIntegerHasher from TColStd); 
							  
    class ListOfCoupleOfShapes  
    	instantiates List from TCollection  (CoupleOfShapes from GEOMAlgo);


    class IndexedDataMapOfShapeState  
    	instantiates IndexedDataMap from TCollection   	(Shape from TopoDS,
	    		    		         	 State from TopAbs,  
	    	    	    	    	    	    	 ShapeMapHasher from TopTools);

end GEOMAlgo;
