--  Copyright (C) 2007-2010  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	GEOMAlgo_ShapeInfoFiller.cdl
--  Created:	Mon Apr  2 15:05:34 2007
--  Author:	Peter KURNEV
--
class ShapeInfoFiller from GEOMAlgo 
    inherits Algo from GEOMAlgo 
     
	---Purpose: 

uses  
    Pln      from gp, 
    Sphere   from gp,
    Cylinder from gp, 
    Cone     from gp, 
    Torus    from gp, 
    
    Shape from TopoDS, 
    Face  from TopoDS,
    Solid from TopoDS, 
     
    ShapeInfo from GEOMAlgo, 
    KindOfName from GEOMAlgo, 
    IndexedDataMapOfShapeShapeInfo from GEOMAlgo

--raises

is  
   
    Create 
    	returns ShapeInfoFiller from GEOMAlgo;   
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_ShapeInfoFiller();"   
    
    SetShape(me:out; 
    	    aS:Shape from TopoDS); 

    Shape(me) 
    	returns Shape from TopoDS; 
    ---C++:return const &  
     
    SetTolerance(me:out; 
    	    aT:Real from Standard);   
	 
    Tolerance(me) 
    	returns Real from Standard;      
     
    Info(me) 
	returns ShapeInfo from GEOMAlgo; 
    ---C++:return const & 

    Info(me; 
    	    aS:Shape from TopoDS) 
	returns ShapeInfo from GEOMAlgo; 
    ---C++:return const & 
     
    Perform(me:out)  
	is redefined;      

    CheckData(me:out) 
	is redefined protected;  
	 
    FillNbSubShapes(me:out; 
    	    aS:Shape from TopoDS; 
    	    aInfo: out ShapeInfo from GEOMAlgo) 
	is protected; 
	 
    FillSubShapes(me:out; 
    	    aS:Shape from TopoDS) 
	is protected; 
	 
    FillShape(me:out; 
    	    aS:Shape from TopoDS) 
	is protected; 
	 
    FillVertex(me:out; 
    	    aS:Shape from TopoDS) 
	is protected; 
     
    FillEdge(me:out; 
    	aS:Shape from TopoDS) 
	is protected; 
  
    FillFace(me:out; 
    	aS:Shape from TopoDS) 
	is protected; 
	 
    FillSolid(me:out; 
    	aS:Shape from TopoDS) 
	is protected; 
     
    FillContainer(me:out; 
    	aS:Shape from TopoDS) 
	is protected; 


    FillDetails(me:out; 
    	    aF:Face from TopoDS; 
    	    aPln:Pln from  gp) 
	is protected; 
	 
    FillDetails(me:out; 
    	    aF:Face from TopoDS; 
    	    aSph:Sphere from gp) 
	is protected;  
     
    FillDetails(me:out; 
    	    aF:Face from TopoDS; 
    	    aCyl:Cylinder from gp) 
	is protected; 
	 
    FillDetails(me:out; 
    	    aF:Face from TopoDS; 
    	    aCone:Cone from gp) 
	is protected;  
	 
    FillDetails(me:out; 
    	    aF:Face from TopoDS; 
    	    aTorus:Torus from gp) 
	is protected;  

    FillDetails(me:out; 
    	    aS:Solid from TopoDS) 
	is protected;    
	
fields
    myShape     : Shape from TopoDS is protected;  
    myEmptyInfo : ShapeInfo from GEOMAlgo is protected;  
    myMapInfo   : IndexedDataMapOfShapeShapeInfo from GEOMAlgo is protected; 
    myTolerance : Real from Standard is protected;
end ShapeInfoFiller;
