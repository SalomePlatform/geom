-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	BlockFix_UnionFaces.cdl
--  Created:	Tue Dec  7 17:15:42 2004
--  Author:	Pavel Durandin
--
class UnionFaces from BlockFix

uses

    Face from TopoDS,
    Shape from TopoDS

is

    Create returns UnionFaces from BlockFix;
    	---Purpose: Empty constructor
    
    GetTolerance(me: in out) returns Real;
    	---Purpose: Returns modifiable tolerance
	---C++: return& 
        
    Perform (me: in out; Shape: Shape from TopoDS) returns Shape from TopoDS;
    	---Purpose: Performs the unification of the fsces
	--          whith the same geometry
	
    IsSameDomain(me; aFace      : Face from TopoDS;
    	    	     aChekedFace: Face from TopoDS)
    returns Boolean is virtual;
    	---Purpose: Returns true is surfaces have same geometrically domain
	--          with given tolerance
	
    MovePCurves(me; aTarget: in out Face from TopoDS;
    	    	    aSource:        Face from TopoDS)
    is virtual;
    	---Purpose: Creates pcurves on aTarget face for each edge from 
	--          aSource one.

fields

    myTolerance: Real;
    
end;
    

