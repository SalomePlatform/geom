--  Copyright (C) 2007-2010  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	NMTTools_CommonBlock.cdl
-- Created:	Tue Dec  9 12:11:48 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class CommonBlock from NMTTools 

	---Purpose: 

uses 
    ListOfInteger   from TColStd, 
    PaveBlock       from BOPTools,
    ListOfPaveBlock from BOPTools

--raises

is 
    Create 
    	returns CommonBlock from NMTTools; 
	 
    AddPaveBlock(me:out; 
	    aPB : PaveBlock from BOPTools); 
	     
    AddFace(me:out; 
	    aF : Integer from Standard); 
	 
    AddFaces(me:out; 
	    aLF:  ListOfInteger from TColStd);    
	     
    PaveBlocks(me) 
    	returns ListOfPaveBlock from BOPTools; 
    ---C++:  return const &  
    
    Faces (me) 
    	returns ListOfInteger from TColStd; 
    ---C++:  return const &  
     
    PaveBlock1  (me) 
    	returns  PaveBlock from BOPTools; 
    ---C++:  return const &	
	 
    PaveBlock1  (me:out; 
    	    anIx: Integer from Standard) 
    	returns  PaveBlock from BOPTools; 
    ---C++:  return & 
     
    PaveBlockOnEdge  (me:out;  
    	    anIndex: Integer from Standard) 
    	returns  PaveBlock from BOPTools; 
    ---C++:  return  &	  
     
    IsPaveBlockOnFace  (me;  
    	    anIndex: Integer from Standard) 
    	returns  Boolean from Standard; 
     
    IsPaveBlockOnEdge  (me;  
    	    anIndex: Integer from Standard) 
    	returns  Boolean from Standard;   
	
    IsEqual  (me; 
    	    aCB:CommonBlock from NMTTools) 
	returns Boolean from Standard; 
	 
    Contains(me; 
    	    aPB:PaveBlock from BOPTools) 
	returns  Boolean from Standard; 
	 
--    SetEdge (me:out;   
--    	    anEdge:Integer from Standard);  

--    Edge (me) 
--    	returns Integer from Standard;  

fields 
    myPaveBlocks: ListOfPaveBlock from BOPTools is protected;  
    myFaces     : ListOfInteger   from TColStd  is protected;  
      	    
end CommonBlock;








