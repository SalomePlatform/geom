-- Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_ShapeSet.cdl
-- Created:	
-- Author:	Peter KURNEV 
--
class ShapeSet from GEOMAlgo 

	---Purpose: Implementation some formal   
    	--          opereations with Set of shapes        

uses 
    Shape from TopoDS,
    MapOfOrientedShape from TopTools, 
    ListOfShape from TopTools,
    ShapeEnum from TopAbs 
    
--raises

is 
    Create 
    	---Purpose: Empty constructor
    	returns ShapeSet from GEOMAlgo; 

    Add(me:out; 
    	    theLS:ListOfShape from TopTools); 
    	---Purpose: Adds shapes from the list theLS to the Set   
	 
    Add(me:out; 
    	    theShape:Shape from TopoDS);
    	---Purpose: Adds shape theShape to the Set 
	
    Add(me:out; 
    	    theShape:Shape from TopoDS; 
    	    theType :ShapeEnum from TopAbs);  
    	---Purpose: Adds sub-shapes of shape theShape, 
    	--          that have type theType to the Set 
	 
    Subtract(me:out; 
	    theSet:ShapeSet from GEOMAlgo); 
    	---Purpose: Removes shapes of theSet from the Set 
	 
    Clear(me:out);
    	---Purpose: Clears internal fields 
	 
    Contains(me; 
	    theSet:ShapeSet from GEOMAlgo) 
    	---Purpose: Returns True if the Set contains  
    	--          all shapes of theSet 
    	returns Boolean from Standard; 
    		     
    GetSet(me) 
    	---Purpose: Returns the Set  
    	returns ListOfShape from TopTools; 
    ---C++: return const &     	 
    --modified by NIZNHY-PKV Wed Oct 28 13:51:45 2010f 
    IsEqual(me; 
	    theOther: ShapeSet from GEOMAlgo) 
    	---Purpose: Returns True if the Set==theSet 
    	returns Boolean from Standard;  
    ---C++: alias operator == 
    --modified by NIZNHY-PKV Wed Oct 28 13:51:50 2010t 
     
fields 
    myMap  : MapOfOrientedShape from TopTools is protected;   
    myList : ListOfShape        from TopTools is protected;

end ShapeSet; 
