-- Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	NMTDS_Iterator.cdl
--  Created:	Sun May 07 14:58:16 2006
--  Author:	Peter KURNEV
--
class Iterator from NMTDS 
     
	---Purpose: 

uses  
    DataMapOfIntegerListOfInteger from TColStd,
    ShapeEnum from TopAbs, 
    ShapesDataStructure  from NMTDS,
    PShapesDataStructure from NMTDS,
    ListOfPassKeyBoolean from NMTDS,
    ListIteratorOfListOfPassKeyBoolean from NMTDS,
    PassKeyBoolean from NMTDS 
    
--raises

is 
    Create   
    	returns Iterator from NMTDS;
    ---C++: alias "Standard_EXPORT virtual ~NMTDS_Iterator();" 
    
   
    SetDS(me:out; 
    	    pDS:PShapesDataStructure from NMTDS); 
     
    DS(me) 
      returns ShapesDataStructure from NMTDS; 
    ---C++:return const & 
     
    Initialize(me: out;  
    	    aType1: ShapeEnum from TopAbs;
    	    aType2: ShapeEnum from TopAbs); 
    More(me)  
    	returns Boolean from Standard; 
  	 
    Next(me: out); 
     
    Current(me; aIndex1:out Integer from Standard;
    	    	aIndex2:out Integer from Standard;
    	    	aWithSubShape: out Boolean from Standard); 
    	
    Prepare(me:out) 
    	is virtual; 
      
    Intersect(me:out) 
    	is virtual protected; 
	
    ExpectedLength(me) 
    	returns Integer from Standard;  
	 
    BlockLength(me) 
    	returns Integer from Standard;  
     
    SDVertices(me) 
    	returns DataMapOfIntegerListOfInteger from TColStd; 
    ---C++:return const &  
     
    FillMVSD(myclass; 
    	aMVSD1:DataMapOfIntegerListOfInteger from TColStd; 
    	aMVSD2:out DataMapOfIntegerListOfInteger from TColStd); 
 
fields
    myDS       :PShapesDataStructure from NMTDS     is protected; 
    myLists    :ListOfPassKeyBoolean from NMTDS [6] is protected;  
    myIterator :ListIteratorOfListOfPassKeyBoolean from NMTDS is protected; 
    myEmptyList:ListOfPassKeyBoolean from NMTDS is protected; 
    myLength   :Integer from Standard is protected; 
    --
    myMVSD     :DataMapOfIntegerListOfInteger from TColStd is protected;     

end Iterator;
