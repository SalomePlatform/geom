// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
// See http://www.salome-platform.org/
//
-- File:	NMTDS.cdl
-- Created:	Fri Nov 28 10:13:19 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2003


package NMTDS 

	---Purpose: 

uses   
    
    TCollection, 
    TColStd,
    Bnd,
    TopoDS, 
    TopAbs, 
    TopTools, 
    BooleanOperations,
    BOPTColStd
is  
    class ShapesDataStructure;
    class IndexRange; 

    pointer PShapesDataStructure to ShapesDataStructure from NMTDS;

    class CArray1OfIndexRange instantiates 
	CArray1 from BOPTColStd(IndexRange from NMTDS); 
     
    class ListOfIndexedDataMapOfShapeAncestorsSuccessors instantiates 
	List from TCollection(IndexedDataMapOfShapeAncestorsSuccessors from BooleanOperations); 
	 
    class IndexedDataMapOfIntegerIndexedDataMapOfShapeInteger instantiates 
    	IndexedDataMap from TCollection(Integer        from Standard, 
	    	    	    	    	IndexedDataMapOfShapeInteger from BooleanOperations, 
					MapIntegerHasher from TColStd); 
					 
end NMTDS;
