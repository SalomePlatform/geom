-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	NMTDS_IteratorCheckerSI.cdl
--  Created:	Tue Feb  6 10:18:27 2007
--  Author:	Peter KURNEV
--
class IteratorCheckerSI from NMTDS  
    inherits Iterator from NMTDS

	---Purpose: 

--uses 
--raises

is 
    Create   
    	returns IteratorCheckerSI from NMTDS;
    ---C++: alias "Standard_EXPORT virtual ~NMTDS_IteratorCheckerSI();" 
     
    Intersect(me:out) 
    	is redefined protected;  
 
--fields
end IteratorCheckerSI;
