-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_Builder.cdl
-- Created:	
-- Author:	Peter KURNEV
--
class Builder from GEOMAlgo 
    	inherits BuilderShape from GEOMAlgo 
	
	---Purpose:   

uses  
    ShapeEnum from TopAbs,
    Shape     from TopoDS, 
     
    ListOfShape                      from TopTools, 
    IndexedDataMapOfShapeListOfShape from TopTools, 
    IndexedDataMapOfShapeShape       from TopTools,   
    MapOfShape                       from TopTools,
    Image     from BRepAlgo, 
    
    PaveFiller from NMTTools, 
    PPaveFiller from NMTTools 
    
--raises

is
 
    Create 
	---Purpose:  Empty constructor     
    	returns Builder from GEOMAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_Builder();" 

    Perform(me:out) 
	---Purpose:  Performs calculations     
    	is redefined; 
	 
    PerformWithFiller(me:out; 
    	theDSF: PaveFiller from NMTTools) 
    	---Purpose:  Performs calculations using prepared PaveFiller 
	--           object theDSF          	 
    	is virtual;
   
    AddShape (me:out;  
    	    theShape: Shape from TopoDS) 
	---Purpose:  Adds argument theShape of the operation    		     
    	is virtual;

    Clear(me:out) 
	---Purpose:  Clears internal fields and arguments             
    	is virtual;  
    
    Shapes(me) 
	---Purpose:  Returns the arguments of the operation       
    	returns ListOfShape from TopTools;  
    ---C++: return const &   
    --
    --  History  support 
    --
    Generated (me:out;  
    	    theS : Shape from TopoDS)
    	---Purpose: Returns the  list of shapes generated from the
    	--          shape theS. 
    	returns ListOfShape from TopTools
    	is redefined;
    	---C++: return const & 

    Modified (me:out;  
    	    theS : Shape from TopoDS)
    	---Purpose: Returns the list of shapes modified from the shape
    	--          theS. 
    	returns ListOfShape from TopTools
    	is redefined;
    	---C++: return const &  

    IsDeleted (me:out;  
    	    theS : Shape from TopoDS) 
    	---Purpose: Returns true if the shape theS has been deleted.
    	returns Boolean from Standard  
    	is redefined; 
    -- 
    --    protected methods  
    --  
    PerformInternal(me:out; 
    	theDSF: PaveFiller from NMTTools) 
    	---Purpose:  Performs calculations using prepared DSFiller 
	--           object theDSF          	 
    	is virtual protected;  
	 
    PrepareHistory (me:out) 
    	---Purpose:  Prepare information for history support  
    	is redefined protected;  
	
    ClearInternals(me:out) 
	---Purpose:  Clears internal fields     
    	is virtual protected;  
      
    Prepare(me:out)  
    	---Purpose:  Provides preparing actions  
    	is virtual protected;   
	 
    PostTreat(me:out)  
    	---Purpose:  Provides post-tratment actions  
    	is virtual protected;
     
    AddShape1 (me:out;  
    	    theShape: Shape from TopoDS) 
    	---Purpose:  Append the argument theShape to  
    	--           typified lists of arguments myShapes1   
    	is protected; 
 
    BuildResult(me:out; 
	    theType: ShapeEnum from TopAbs) 
    	---Purpose: Build the resulting shapes of type theType      
    	is virtual protected;  
	
    --  Vertices 
    FillImagesVertices(me:out)  
    	---Purpose: Fill Images for vertices   
    	is protected; 
	 
    --  Edges 
    FillImagesEdges(me:out) 
    	---Purpose: Fill Images for edges  
    	is protected; 
    -- 
    --  Faces 
    FillImagesFaces(me:out)  
    	---Purpose: Fill Images for faces 
    	is protected; 
 
    FillIn2DParts(me:out)  
    	---Purpose: For each interferred face find split edges 
	--          that are in 2-D domain of the face           
    	is protected; 
	  
    BuildSplitFaces(me:out)  
    	---Purpose: Build draft faces    
    	is protected; 
	 
    FillSameDomainFaces(me:out)  
    	---Purpose: Among draft faces find same domain faces 
    	is protected; 
 
    FillImagesFaces1(me:out) 
    	---Purpose: Fill Images for faces  
        --          taking into account same domain faces   	 
    	is protected;  
	
    FillInternalVertices(me:out)  
    	---Purpose: Update Images for faces by  
    	--          internal vertices    
    	is protected;  
    -- 
    --  Wires, Shells, Compsolids, Compounds
    FillImagesContainers(me:out; 
    	    theType:ShapeEnum from TopAbs) 
	---Purpose:  Fill Images for Wires, Shells, Compsolids, Compounds        
    	is protected;   
    -- 
    --  Solids  
    FillImagesSolids(me:out)  
    	---Purpose:  Fill Images for solids
    	is protected;  
    	 
    FillIn3DParts(me:out) 
    	---Purpose: For each interferred solid find split faces 
	--          that are in 3-D domain of the solid   
    	is protected; 
 
    BuildSplitSolids(me:out) 
    	---Purpose: Build draft solids   
    	is protected; 
	 
    FillInternalShapes(me:out)  
    	---Purpose:  Update draft solids by 
	--           internal shells, edges, vertices 				     
    	is protected;  
	 
    BuildDraftSolid(me:out; 
    	    theSolid: Shape from TopoDS; 
    	    theDraftSolid: out Shape from TopoDS; 
    	    theInternalFaces: out ListOfShape from TopTools)  
    	---Purpose:  Build solid theDraftSolid that consists of  
    	--           non-internal split faces of the solid   
        --           theSolid.  
    	--           All splits of internal faces of 
        --           theSolid are in the list: theInternalFaces    	 
    	is protected;   
    -- 
    --  debug  methods  
    --
    AddCompound (me:out;  
    	    theShape: Shape from TopoDS); 
	---Purpose:  Adds arguments of the operation as  
        --           shapes of upper level of container shape theShape    	  
    Shapes1(me; 
    	    theType: Integer from Standard) 
        ---Purpose: Returns list of arguments of type theType      	     
    	returns ListOfShape from TopTools; 
    ---C++: return const & 
     
    Images(me)  
    	---Purpose: Returns image shapes    
    	returns Image from BRepAlgo; 
    ---C++: return const &  

    InParts(me; 
    	    theShape:Shape from TopoDS)  
	---Purpose: Returns split-parts of shapes that have  
        --          state IN for the domain of shape theShape    	 
    	returns ListOfShape from TopTools; 
    ---C++: return const &  
 
    -- =====================================================
 
fields 
    myPaveFiller      : PPaveFiller from NMTTools is protected;  
    myShapes          : ListOfShape from TopTools is protected; 
    -- Common usage 
    myNbTypes         : Integer from Standard is protected; 
    myMapFence        : MapOfShape from TopTools is protected;        
    myShapes1         : ListOfShape from TopTools[9] is protected; 
    myImages          : Image from BRepAlgo is protected;  
    myInParts         : IndexedDataMapOfShapeListOfShape from TopTools is protected; 
     
    -- Faces
    mySplitFaces      : Image from BRepAlgo is protected;  
    mySameDomainShapes: IndexedDataMapOfShapeShape from TopTools is protected;
    --  solids 
    myDraftSolids     : IndexedDataMapOfShapeShape from TopTools is protected; 
    myEntryPoint      : Integer from Standard is protected;
    --     
end Builder;

