--  GEOM PARTITION : partition algorithm
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : Partition_Spliter.cdl
--  Author : Benedicte MARTIN
--  Module : GEOM

class Spliter from Partition

        ---Purpose: Split solids, shells and  faces  into parts of the
        --          same  topology  if  reconstruction  level  is  not
        --          limited.

uses
    Inter3d             from Partition,
    Loop2d              from Partition,
    Builder             from BRep,
    ShapeEnum           from TopAbs,
    Compound            from TopoDS,
    Face                from TopoDS,
    Edge                from TopoDS,
    Shape               from TopoDS,
    MapOfOrientedShape  from TopTools,
    IndexedMapOfShape   from TopTools,
    DataMapOfShapeShape from TopTools,
    ListOfShape         from TopTools,
    MapOfShape          from TopTools,
    AsDes               from BRepAlgo,
    Image               from BRepAlgo

is
    Create  returns Spliter from Partition;
        ---Purpose: constructor

    AddShape ( me : in out; S : Shape from TopoDS);
        ---Purpose: add object Shape to be splitted.
        --          If S  is  a  COMPOUND  or  COMPSOLID,  it  will be
        --          exploded  in  order  to  get  more  simple  object
        --          shapes. 
        --          Object shapes that  are  vertices,  edges or wires
        --          won't be splitted and won't be in a result.

    AddTool  ( me : in out; S : Shape from TopoDS);
        ---Purpose: add cutting tool

    Compute (me : in out; Limit : ShapeEnum from TopAbs
                          = TopAbs_SHAPE);
        ---Purpose: produce a result which  is  a compound of parts of
        --          object shapes.  A  part  can  be  either a vertex,
        --          edge, wire, face, shell or solid.
        --          By default, a part is  of  the same topology as an
        --          object  shape,   else   <Limit>   restricts  parts
        --          reconstruction.
        --          If <Limit> == TopAbs_VERTEX, only new vertices are
        --          returned in the result

    KeepShapesInside (me : in out; S : Shape from TopoDS);
        ---Purpose: remove shapes that are outside of S from result.
        --          S should be an object shape.
        ---Warning: call it after Compute()

    RemoveShapesInside (me : in out; S : Shape from TopoDS);
        ---Purpose: remove shapes that are inside S from result.
        --          S should be an object shape.
        ---Warning: call it after Compute()

    Shape ( me ) returns Shape from TopoDS;
        ---Purpose: return resulting compound

    Clear ( me : in out);
        ---Purpose: clear fields


        ---Category: private methods


    MakeSolids (me: in out; Solid : Shape from TopoDS;
                            Shells: in out ListOfShape from TopTools) 
        is private;
        ---Purpose: make solids out of Shells

    MakeShells (me: in out; S : Shape from TopoDS;
                            NS: in out ListOfShape from TopTools) is private;
        ---Purpose: split S into shells

    MakeFaces (me: in out; S : Shape from TopoDS)
        returns Shape from TopoDS is private;
        ---Purpose: split faces of S, return compound of new faces

    MakeEdges (me; 
               E : Edge from TopoDS;
               VOnE : ListOfShape from TopTools;
               NE : in out ListOfShape from TopTools) 
        is private;
        ---Purpose: cut E by vertices  VOnE,  return list of new edges
        --          NE
    
    FindFacesInside (me: in out; S : Shape from TopoDS;
                                 CheckClosed : Boolean = Standard_False;
                                 All         : Boolean = Standard_False)
        returns Shape from TopoDS is private;
        ---Purpose: return compound of faces  of other shapes that are
        --          inside <S>. <S>  must  have image in myImageShape.
        --          <CheckClosed> makes avoid faces that do not form a
        --          closed shell
        --          <All> makes return already added faces

    CheckTool ( me: in out; S : Shape from TopoDS)
        returns Boolean from Standard is private;
        ---Purpose: Return True if <S>  is  a tool shape. Prepare tool
        --          faces of <S> for the search of internal faces.

    MergeEqualEdges (me: in out; LE : ListOfShape from TopTools) is private;
        ---Purpose: among LE, find  equal  edges,  choose ones to keep
        --          and make them have  pcurves  on all faces they are
        --          shared by
        --          <LE> contains edge splits

    IsInside (myclass; S1,S2 : Shape from TopoDS)
        returns Boolean from Standard is private;
        ---Purpose: Return True if the first vertex of S1 inside S2.
        --          If S1.IsNull(), check infinite point against S2.

    GetOriginalShape(me; aShape : Shape from TopoDS)
        returns Shape from TopoDS is private;
        ---Purpose: Return the  shape  aShape  originates from. aShape
        --          should be a face or more complex result shape

    FindToolsToReconstruct(me: in out) is private;
        ---Purpose: find and store  as  objects  tools which interfere
        --          with  solids   or   are   inside   solids  without
        --          an interference

fields

    myDoneStep     : ShapeEnum           from TopAbs;   -- rebuilt level
    myShape        : Compound            from TopoDS;   -- result
    myBuilder      : Builder             from BRep;
    		   			   
    myListShapes   : ListOfShape         from TopTools; -- object shapes
    myMapFaces     : MapOfShape          from TopTools; -- object faces
    myMapTools     : MapOfShape          from TopTools; -- tool faces
    myEqualEdges   : MapOfShape          from TopTools; -- equal splits
    myNewSection   : MapOfShape          from TopTools; -- new secton edges
    myClosedShapes : MapOfShape          from TopTools;
    myWrappingSolid: MapOfShape          from TopTools; -- solids having other shapes inside
    myFaceShapeMap : DataMapOfShapeShape from TopTools; -- to find a shape by face
    		   			   
    myInternalFaces: DataMapOfShapeShape from TopTools; -- shape and its internal faces
    myIntNotClFaces: DataMapOfShapeShape from TopTools; -- internal but not closed 

		   			   
    myAsDes        : AsDes               from BRepAlgo;
    myImagesFaces  : Image               from BRepAlgo;   
    myImagesEdges  : Image               from BRepAlgo;    
    myImageShape   : Image               from BRepAlgo;
    
        -- contains info of same domain shapes and section edges
    myInter3d      : Inter3d             from Partition;
    
        -- avoid rebuilding twice commont part of solids
    myAddedFacesMap: MapOfOrientedShape  from TopTools;
    
end Spliter;
