-- Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	NMTTools_Tools.cdl
-- Created:	Mon Dec  8 10:32:34 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class Tools from NMTTools 

	---Purpose: 

uses
    Vertex from TopoDS, 
    Edge from TopoDS, 
    Face from TopoDS, 
    Context from IntTools,  
    Curve from Geom2d,
     
    ListOfShape from TopTools,
    IndexedDataMapOfIntegerIndexedMapOfInteger from BOPTColStd, 
    CArray1OfVVInterference from BOPTools, 
    CArray1OfSSInterference from BOPTools, 
    ListOfCoupleOfShape from NMTTools, 
    IndexedDataMapOfShapeIndexedMapOfShape from NMTTools

--raises

is 
    MakeNewVertex  (myclass;  
        	    aLV : ListOfShape from TopTools; 
		    aNewVertex: out Vertex from TopoDS); 
    FindChains(myclass; 
    	aVVs:CArray1OfVVInterference from BOPTools; 
	aMCX: out IndexedDataMapOfIntegerIndexedMapOfInteger from BOPTColStd); 
     
    FindChains(myclass; 
    	aVVs:CArray1OfSSInterference from BOPTools; 
	aMCX: out IndexedDataMapOfIntegerIndexedMapOfInteger from BOPTColStd);  
     
    FindChains(myclass;   
    	aMCV: IndexedDataMapOfIntegerIndexedMapOfInteger from BOPTColStd; 
	aMCX: out IndexedDataMapOfIntegerIndexedMapOfInteger from BOPTColStd); 
	
     
    IsSplitInOnFace(myclass; 
    	    aE  : Edge from TopoDS; 
	    aF  : Face from TopoDS; 
	    aCtx: Context from IntTools) 
    	returns Boolean from Standard; 

    AreFacesSameDomain(myclass; 
	    aF1  : Face from TopoDS; 
	    aF2  : Face from TopoDS; 
    	    aCtx : Context from IntTools) 
    	returns Boolean from Standard; 

    FindChains(myclass; 
    	    aLCS:ListOfCoupleOfShape from NMTTools; 
	    aM  :out  IndexedDataMapOfShapeIndexedMapOfShape from NMTTools);	

    FindChains(myclass; 
    	    aM1: IndexedDataMapOfShapeIndexedMapOfShape from NMTTools;
	    aM2:out  IndexedDataMapOfShapeIndexedMapOfShape from NMTTools);

    MakePCurve(myclass;  
    	    aE   :  Edge from TopoDS; 
    	    aF   :  Face from TopoDS;  
    	    aC2D :  Curve from Geom2d); 
	     
    UpdateEdge(myclass;  
    	    aE   :  Edge from TopoDS;   
    	    aTol :  Real from Standard);	
--fields

end Tools;
