-- File:	NMTTools_CommonBlock.cdl
-- Created:	Tue Dec  9 12:11:48 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2003


class CommonBlock from NMTTools 

	---Purpose: 

uses 
    ListOfInteger   from TColStd, 
    PaveBlock       from BOPTools,
    ListOfPaveBlock from BOPTools

--raises

is 
    Create 
    	returns CommonBlock from NMTTools; 
	 
    AddPaveBlock(me:out; 
	    aPB : PaveBlock from BOPTools); 
	     
    AddFace(me:out; 
	    aF : Integer from Standard); 
	 
    AddFaces(me:out; 
	    aLF:  ListOfInteger from TColStd);    
	     
    PaveBlocks(me) 
    	returns ListOfPaveBlock from BOPTools; 
    ---C++:  return const &  
    
    Faces (me) 
    	returns ListOfInteger from TColStd; 
    ---C++:  return const &  
     
    PaveBlock1  (me) 
    	returns  PaveBlock from BOPTools; 
    ---C++:  return const &	
	 
    PaveBlock1  (me:out; 
    	    anIx: Integer from Standard) 
    	returns  PaveBlock from BOPTools; 
    ---C++:  return & 
     
    PaveBlockOnEdge  (me:out;  
    	    anIndex: Integer from Standard) 
    	returns  PaveBlock from BOPTools; 
    ---C++:  return  &	  
     
    IsPaveBlockOnFace  (me;  
    	    anIndex: Integer from Standard) 
    	returns  Boolean from Standard; 
     
    IsPaveBlockOnEdge  (me;  
    	    anIndex: Integer from Standard) 
    	returns  Boolean from Standard;   
	
    IsEqual  (me; 
    	    aCB:CommonBlock from NMTTools) 
	returns Boolean from Standard; 
	 
    Contains(me; 
    	    aPB:PaveBlock from BOPTools) 
	returns  Boolean from Standard; 
	 
--    SetEdge (me:out;   
--    	    anEdge:Integer from Standard);  

--    Edge (me) 
--    	returns Integer from Standard;  

fields 
    myPaveBlocks: ListOfPaveBlock from BOPTools is protected;  
    myFaces     : ListOfInteger   from TColStd  is protected;  
      	    
end CommonBlock;








