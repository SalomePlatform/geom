--  Copyright (C) 2007-2010  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_Gluer1.cdl
-- Created:	Wed Jan 24 11:37:31 2007
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class Gluer1 from GEOMAlgo  
    inherits  Gluer from GEOMAlgo

	---Purpose: 

uses 
    ListOfCoupleOfShapes from GEOMAlgo, 
    DataMapOfPassKeyShapeShape from GEOMAlgo 

--raises

is 
    Create   
    	returns Gluer1 from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_Gluer1();" 
      
    SetFacesToUnglue(me:out; 
    	aLCS:ListOfCoupleOfShapes from GEOMAlgo);
	 
    FacesToUnglue(me) 
    	returns ListOfCoupleOfShapes from GEOMAlgo;  	        	
    ---C++: return const& 
       
    GluedFaces(me) 
    	returns ListOfCoupleOfShapes from GEOMAlgo;  	        	
    ---C++: return const&  
      
    RejectedFaces(me) 
    	returns ListOfCoupleOfShapes from GEOMAlgo;  	        	
    ---C++: return const&   
    
    Perform(me:out) 
	is redefined; 
     
    UnglueFaces(me:out); 
     
    FillGluedFaces(me:out) 
     	is protected; 
	
fields
    myGluedFaces        :ListOfCoupleOfShapes from GEOMAlgo is protected;
    myFacesToUnglue     :ListOfCoupleOfShapes from GEOMAlgo is protected;
    myRejectedFaces     :ListOfCoupleOfShapes from GEOMAlgo is protected; 
    myMapGN             :DataMapOfPassKeyShapeShape from GEOMAlgo is protected; 

end Gluer1;
