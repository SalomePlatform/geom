--  Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

--  File:	GEOMAlgo_ShapeAlgo.cdl
--  Created:	Tue Dec  7 12:05:19 2004
--  Author:	Peter KURNEV
--
deferred class ShapeAlgo from GEOMAlgo 
    inherits Algo from GEOMAlgo  
    
	---Purpose: 

uses
    Shape from TopoDS, 
    Context from IntTools

--raises

is
    Initialize 
    	returns ShapeAlgo from GEOMAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_ShapeAlgo();"  
    
    SetShape(me:out; 
    	    aS:Shape from TopoDS);
     
    SetTolerance(me:out; 
    	    aT:Real from Standard); 
	     
    Shape(me) 
    	returns Shape from TopoDS; 
    ---C++:return const &  
     
    Tolerance(me) 
    	returns Real from Standard;  
     
    Result(me) 
    	returns Shape from TopoDS; 
    ---C++:return const &  
    
fields 
    myShape     : Shape from TopoDS is protected;     
    myTolerance : Real from Standard is protected; 
    myResult    : Shape from TopoDS is protected; 
    myContext   : Context from IntTools is protected; 
    
end ShapeAlgo;
