-- File:	GEOMAlgo_VertexSolid.cdl
-- Created:	Wed Jan 12 16:34:53 2005
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2005


class VertexSolid from GEOMAlgo  
    	inherits ShapeSolid from GEOMAlgo

	---Purpose: 

--uses
--raises

is
    Create   
    	returns  VertexSolid from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_VertexSolid();"
     
    Perform (me:out) 
	is redefined; 
	 
    Prepare(me:out)  
   	 is redefined protected;
     
    BuildResult (me:out) 
	is redefined protected; 
    
--fields

end VertexSolid;
