-- File:	GEOMAlgo_PassKey.cdl
-- Created:	
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 


class PassKey from GEOMAlgo 

	---Purpose: 

uses
    Shape from TopoDS, 
    ListOfInteger from TColStd   
  	 
--raises

is 
    Create  
    	returns PassKey from GEOMAlgo; 
     
    Assign(me:out;  
    	    Other : PassKey from GEOMAlgo) 
    	returns PassKey from GEOMAlgo; 
    ---C++: alias operator =
    ---C++: return & 
--    
    SetIds(me:out; 
    	    aI1  :Integer from Standard); 
	     
    SetIds(me:out; 
    	    aI1 :Integer from Standard;    
    	    aI2 :Integer from Standard);  
	     
    SetIds(me:out; 
    	    aI1 :Integer from Standard;    
    	    aI2 :Integer from Standard;    
    	    aI3 :Integer from Standard);  

    SetIds(me:out; 
    	    aI1 :Integer from Standard;    
    	    aI2 :Integer from Standard;    
    	    aI3 :Integer from Standard;    
    	    aI4 :Integer from Standard); 
     
    SetIds(me:out;  
    	    aLS  :ListOfInteger from TColStd);   
 
    NbMax(me) 
	returns Integer  from Standard; 
	 
    Clear(me:out); 
     
    Compute(me:out); 
     
    IsEqual(me; 
    	    aOther:PassKey from GEOMAlgo) 
	returns Boolean from Standard;   		     

    Key(me) 
    	returns Address from Standard;  
	 
    HashCode(me; 
	    Upper : Integer  from Standard)  
    	returns Integer from Standard;   	 
     
    Id(me; 
    	    aIndex: Integer  from Standard)  
    	returns Integer from Standard;
    	

    Dump(me); 

fields 
 
    myNbIds: Integer from Standard is protected;  
    myNbMax: Integer from Standard is protected; 
    mySum  : Integer from Standard is protected;   
    myIds  : Integer from Standard [8] is protected; 

end PassKey;
