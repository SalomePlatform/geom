-- File   :	Partition_Loop2d.cdl
-- Created:	Thu Aug 02 16:07:39 2001
-- Author :	Benedicte MARTIN
--		
---Copyright:	 OPEN CASCADE 2001


class Loop2d from Partition

        ---Purpose: Builds the loops from a set of edges on a face.
	--          It works in  supposition  that  all constant edges
	--          are split edges of  an initialization face and all
	--          section edges are new on the face

uses

    Orientation               from TopAbs,
    Boolean                   from Standard,
    Face                      from TopoDS,
    Image                     from BRepAlgo,
    Face                      from TopoDS,
    Edge                      from TopoDS,
    ListOfShape               from TopTools,
    DataMapOfShapeListOfShape from TopTools,
    MapOfShape                from TopTools
is

    Create;
    
    Init (me : in out; F : Face from TopoDS)
	---Purpose: Init with <F> the set of edges must have
	--          pcurves on <F>. 
    is static;
    
    AddConstEdge  (me : in out; E : Edge from TopoDS)
	---Purpose: Add <E> as unique edge in the result.
    is static;

    AddSectionEdge  (me : in out; E : Edge from TopoDS)
	---Purpose: Add <E> as double edge in the result.
    is static;

    Perform(me : in out)
	---Purpose: Make loops.
    is static;
    
    NewWires (me)	
	---Purpose: Returns the list of wires performed. 
	--          can be an empty list.
	---C++: return const &
    returns ListOfShape from TopTools;
    	
    WiresToFaces (me : in out; EdgeImage : Image      from BRepAlgo)
    	---Purpose:  Build faces from the wires result.
    	--           <EdgeImage> serves to  find  original edge by new
    	--           one.
    is static;
    
    NewFaces (me)
        ---Purpose: Returns the list of faces.
    	---Warning: The method <WiresToFaces> as to be called before.
    	--          can be an empty list.
	---C++: return const &
    returns ListOfShape from TopTools;

    
fields

    myFace       : Face        from TopoDS;
    myFaceOri    : Orientation from TopAbs;
    myConstEdges : ListOfShape from TopTools;
    myNewWires   : ListOfShape from TopTools;
    myNewFaces   : ListOfShape from TopTools;

     -- internal wires do not contain constant edges
    myInternalWL : ListOfShape from TopTools;
    
    mySectionEdges : MapOfShape from TopTools;
    
end Loop2d;
