-- File:	GEOMAlgo_SolidSolid.cdl
-- Created:	Wed Jan 26 12:05:14 2005
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2005


class SolidSolid from GEOMAlgo 
    inherits ShellSolid from GEOMAlgo 
    
	---Purpose: 

uses 
    Shape from TopoDS

--raises

is
    Create   
    	returns SolidSolid from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_SolidSolid();" 
    
    Perform (me:out) 
	is redefined; 
	 
    BuildResult (me:out) 
	is redefined protected; 	
    
    SetShape2 (me:out;  
    	    aS: Shape from TopoDS);

    Shape2 (me)  
    	returns Shape from TopoDS; 
    ---C++: return const &  

fields
    myS2: Shape from TopoDS is protected; 
    
end SolidSolid;
