// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
//
-- File:	NMTAlgo_Algo.cdl
-- Created:	Tue Jan 27 14:41:04 2004
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2004


deferred class Algo from NMTAlgo 

	---Purpose: 

uses 
    Shape     from TopoDS, 
    
    DSFiller  from NMTTools,
    PDSFiller from NMTTools

--raises

is
    Initialize 
    	returns Algo from NMTAlgo;  
    ---C++: alias "Standard_EXPORT virtual ~NMTAlgo_Algo();" 
      
     
    SetFiller(me:out; 
    	    aDSF: DSFiller from NMTTools);
     
    Filler(me)
    	returns DSFiller from NMTTools; 
    ---C++:  return const &     
     
    ComputeWithFiller(me:out; 
    	aDSF: DSFiller from NMTTools) 
    	is virtual;  
	 
    Clear (me:out) 
    	is virtual; 
	
    Shape (me) 
     	returns Shape from TopoDS;
    ---C++:  return const &  	 	    		  
     
    IsDone(me) 
    	returns Boolean from Standard; 
     
    ErrorStatus (me) 
    	returns Integer from Standard; 

fields 
    myDSFiller       : PDSFiller from NMTTools   	is protected; 
    myShape          : Shape   from TopoDS      	is protected;
    -- 
    myIsDone         : Boolean from Standard    	is protected; 
    myIsComputed     : Boolean from Standard    	is protected; 
    myErrorStatus    : Integer from Standard    	is protected;	 
    myDraw           : Integer from Standard   	        is protected;  
    
end Algo;
