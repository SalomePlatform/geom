-- File:	GEOMAlgo_FinderShapeOn.cdl
-- Created:	Tue Jan 11 14:35:52 2005
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2005


class FinderShapeOn from GEOMAlgo 
    inherits ShapeAlgo from GEOMAlgo 
    
	---Purpose: 

uses
    Surface from Geom, 
    ShapeEnum from TopAbs, 
    ListOfShape from TopTools, 
    DataMapOfShapeShape from TopTools, 
    Shape from TopoDS, 
    State from GEOMAlgo, 
    IndexedDataMapOfShapeState from GEOMAlgo 
    
--raises

is 
    Create   
    	returns FinderShapeOn from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_FinderShapeOn();" 
     
    Perform(me:out) 
	is redefined;  
	 
    SetSurface(me:out; 
    	    aS:Surface from Geom); 
	 
    SetShapeType(me:out; 
    	    aST:ShapeEnum from TopAbs); 
	 
    SetState(me:out; 
    	    aSF:State from GEOMAlgo);      
     
    Surface(me) 
    	returns Surface from Geom; 
    ---C++: return const & 
     
    ShapeType(me) 
    	returns ShapeEnum from TopAbs; 
	 
    State(me)
    	returns State from GEOMAlgo;  
     
    Shapes(me)
	returns ListOfShape from TopTools; 
    ---C++: return const &  
     
    -- 
    --  protected  methods
    -- 
    CheckData(me:out) 
	is redefined protected; 

    MakeArgument1(me:out) 
	is protected;  

    MakeArgument2(me:out) 
	is protected;
     
    Find(me:out) 
	is protected; 

    Find(me:out; 
    	    aS:Shape from TopoDS) 
	is protected; 

    FindVertices(me:out) 
	is protected; 
	 
    CopySource(myclass; 
    	aS  :Shape from TopoDS; 
	aImages   : out DataMapOfShapeShape from TopTools;   	 
	aOriginals: out DataMapOfShapeShape from TopTools;   	 
    	aSC : out Shape from TopoDS); 
	
					

fields 
    mySurface    : Surface from Geom is protected;  
    myShapeType  : ShapeEnum from TopAbs is protected;  
    myState      : State from GEOMAlgo is protected; 
    myArg1       : Shape from TopoDS is protected;  
    myArg2       : Shape from TopoDS is protected;  
    myLS         : ListOfShape from TopTools is protected;
    myImages     : DataMapOfShapeShape from TopTools is protected; 
    myMSS        : IndexedDataMapOfShapeState from GEOMAlgo is protected; 
    myIsAnalytic : Boolean from Standard is protected; 
     
end FinderShapeOn;
