--  Copyright (C) 2007-2010  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_WireEdgeSet.cdl
-- Created:	
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class WireEdgeSet from GEOMAlgo 

	---Purpose: 

uses
    Face   from TopoDS, 
    Shape  from TopoDS, 
    ListOfShape from TopTools
--raises

is 
    Create   
    	returns WireEdgeSet from GEOMAlgo;  
	 
    Clear(me:out);
	 
    SetFace(me:out; 
    	    aF:Face from TopoDS); 
	     
    Face(me) 
	 returns Face from TopoDS; 
    ---C++: return const &  
     
    AddStartElement(me:out; 
    	    sS: Shape from TopoDS);  
	    
    StartElements(me)  
    	returns ListOfShape from TopTools;
    ---C++: return const & 

    AddShape(me:out; 
    	    sS:Shape from TopoDS); 
	     
    Shapes(me)  
    	returns ListOfShape from TopTools;
    ---C++: return const & 

fields
    myFace         : Face from TopoDS is protected; 
    myStartShapes  : ListOfShape from TopTools is protected;
    myShapes       : ListOfShape from TopTools is protected;  
    
end WireEdgeSet;
