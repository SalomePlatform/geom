-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	NMTTools_CoupleOfShape.cdl
-- Created:	Wed Jan 28 15:03:39 2004
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class CoupleOfShape from NMTTools 

	---Purpose: 

uses
    Shape from TopoDS 
    
--raises

is 
    Create 
    	returns CoupleOfShape from NMTTools; 

    SetShape1(me:out; 
    	aS: Shape from TopoDS); 
	 
    SetShape2(me:out; 
    	aS: Shape from TopoDS); 
	 
    Shape1(me) 
    	returns Shape from TopoDS; 
    ---C++: return const & 	 

    Shape2(me) 
    	returns Shape from TopoDS; 
    ---C++: return const & 
    
fields 
    myShape1:Shape from TopoDS is protected;    
    myShape2:Shape from TopoDS is protected;    

end CoupleOfShape;
