// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
//
-- File:	BlockFix_UnionEdges.cdl
-- Created:	Tue Dec  7 15:24:51 2004
-- Author:	Sergey KUUL
--		<skl@novgorox.nnov.matra-dtv.fr>

class UnionEdges from BlockFix

    	---Purpose: 
	
uses
    
    Shape           from TopoDS,
    ReShape         from ShapeBuild

is

    Create returns UnionEdges from BlockFix;
    
    Perform(me: in out; Shape: Shape from TopoDS;
                        Tol  : Real)
    returns Shape from TopoDS;    
    
fields

    myTolerance : Real;
    myContext   : ReShape from ShapeBuild;
    
end UnionEdges;
