-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_ClsfSurf.cdl
-- Created:	Wed Nov 22 10:19:29 2006
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
class ClsfSurf from GEOMAlgo 
    inherits Clsf from GEOMAlgo 
     
	---Purpose: 

uses  
    Curve   from Geom, 
    Surface from Geom,
    Surface from GeomAdaptor 
    
--raises

is 
    Create 
    	returns mutable ClsfSurf from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_ClsfSurf();"  
      
    SetSurface(me:mutable; 
    	    aS:Surface from Geom);  
	 
    Surface(me) 
    	returns Surface from Geom; 
    ---C++: return const &     
     
    Perform(me:mutable) 
	is redefined;      

    CheckData(me:mutable) 
	is redefined;  
    	
    CanBeON(me; 
    	    aC:Curve from Geom) 
	returns Boolean from Standard 
    	is redefined; 

    CanBeON(me; 
    	    aST:Surface from Geom) 
	returns Boolean from Standard 
    	is redefined;   
	 
fields 
    myS   : Surface from Geom is protected;   
    myGAS : Surface from GeomAdaptor is protected; 
    
end ClsfSurf;
