-- File:	NMTTools_PaveFiller.cdl
-- Created:	Fri Dec  5 14:35:00 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2003


class PaveFiller from NMTTools 

	---Purpose: 

uses    
    ListOfInteger from TColStd,
    Pnt from gp,
    ShapeEnum  from  TopAbs, 
    Vertex     from  TopoDS, 
    Face       from  TopoDS, 
    
    Context     from IntTools, 
    ShrunkRange from IntTools,
      
    IndexedDataMapOfShapeInteger from BooleanOperations, 
    
    InterferencePool  from BOPTools,
    PInterferencePool from BOPTools, 
    PavePool          from BOPTools, 
    PaveBlock         from BOPTools,
    ListOfPaveBlock   from BOPTools,
    SplitShapesPool   from BOPTools, 
    Pave              from BOPTools, 
    PaveSet           from BOPTools, 
    Curve             from BOPTools, 
    SSInterference    from BOPTools, 
    
    IDMapOfPaveBlockIMapOfPaveBlock from BOPTools, 
    IDMapOfPaveBlockIMapOfInteger   from BOPTools, 
    SSIntersectionAttribute         from BOPTools, 
    
    CommonBlockPool         from NMTTools, 
    CommonBlock             from NMTTools, 
    ListOfCommonBlock       from NMTTools,
    IteratorOfCoupleOfShape from NMTTools,
    
    ShapesDataStructure  from NMTDS, 
    PShapesDataStructure from NMTDS 
    
--raises

is 
    Create 
    	returns PaveFiller from NMTTools; 
      
    Create(aIP:InterferencePool from BOPTools)
    	returns PaveFiller from NMTTools; 
     
    Destroy (me: in out) 
	is  virtual;    
    ---C++: alias "Standard_EXPORT virtual ~NMTTools_PaveFiller(){Destroy();}"
    -- 
    --  Selectors/Modifiers
    SetInterferencePool(me:out; 
    	    aIP:InterferencePool from BOPTools);
    
    InterfPool(me:out) 
    	returns PInterferencePool from BOPTools; 
    --	 
    --  Perform the algo  
    Init       (me:out) 
	is protected; 
	 
    Perform    (me:out) 
	is virtual;   
	 
    PerformVV  (me:out) 
    	is virtual protected;  
     
    PerformVE  (me:out) 
    	is virtual protected; 
     
    PerformVF  (me:out) 
    	is virtual protected; 

    PerformEE (me:out) 
    	is virtual protected; 
      
    PerformEF (me:out) 
    	is virtual protected; 
   
    PerformFF (me:out) 
    	is virtual protected; 
     
    MakeSplitEdges(me:out) 
    	is protected;   
     
    PreparePaveBlocks (me:out; 
    	    aType1: ShapeEnum  from  TopAbs; 
    	    aType2: ShapeEnum  from  TopAbs) 
    	is virtual protected; 
     
    CorrectShrunkRanges(me:out; 
    	    aSide:  Integer  from  Standard; 
    	    aPave:  Pave from BOPTools; 
    	    aSR  :  out ShrunkRange  from  IntTools)
    	is protected; 
	 
    PreparePaveBlocks (me:out;   
    	    anE:Integer from Standard) 
    	is virtual protected;  		  
		       
    PerformNewVertices  (me:out) 
    	is virtual protected;  
     
    PrepareEdges  (me:out) 
    	is virtual protected;  
     
    SortTypes      (me;   
    	    anInd1:in out Integer from Standard; 
            anInd2:in out Integer from Standard) 
    	is protected; 
     
    ExpectedPoolLength(me) 
    	returns  Integer from Standard 
	is protected;  
    --
    -- Query section 
    IsDone(me) 
    	returns  Boolean from Standard; 

    DS(me:out) 
    	returns PShapesDataStructure from NMTDS;  
	 
    Context(me) 
    	 returns Context from IntTools; 
    	---C++:return const &	

    ChangeContext(me:out) 
    	 returns Context from IntTools;  
    	---C++:return &	

    PavePool(me) 
    	returns  PavePool from BOPTools; 
    	---C++:return const &	 

    ChangePavePool(me:out) 
    	returns  PavePool from BOPTools; 
    	---C++:return &	

    CommonBlockPool(me) 
    	returns  CommonBlockPool from NMTTools; 
    	---C++:return const &	 

    ChangeCommonBlockPool(me:out) 
    	returns  CommonBlockPool from NMTTools; 
    	---C++:return &	

    SplitShapesPool(me)  
    	returns  SplitShapesPool from BOPTools;
    	---C++:return const &	

    ChangeSplitShapesPool(me:out)  
    	returns  SplitShapesPool from BOPTools;
    	---C++:return  &	
     
    FindSDVertex (me; 
    	    	    nV:  Integer  from  Standard) 
    	returns Integer from Standard; 

    IsSuccesstorsComputed (me;  
    	    iF1:Integer from  Standard; 
    	    iF2:Integer from  Standard) 
    	returns  Boolean from Standard 
    	is protected;  

    IsBlocksCoinside (me; 
    	    aPB1:PaveBlock from BOPTools;
    	    aPB2:PaveBlock from BOPTools) 
	returns Boolean from Standard 
    	is protected; 
     
    RefinePavePool(me:out) 
    	is protected;  

    CheckFacePaves(me:out;  
    	     aV : Vertex  from TopoDS;  
     	     nF:  Integer from Standard) 
    	returns Integer from Standard 
    	is protected;  
	 
    ReplaceCommonBlocks (me:out; 
	    aLCB: ListOfCommonBlock from NMTTools) 
        is protected; 
     
    RemoveCommonBlocks (me:out; 
	    aLCB: ListOfCommonBlock from NMTTools) 
        is protected;
     
    SplitCommonBlocks (me:out; 
	    aLCB: ListOfCommonBlock from NMTTools) 
        is protected;  

    SplitCommonBlock (me:out; 
    	    aCB : CommonBlock from NMTTools; 
	    aLCB: out ListOfCommonBlock from NMTTools) 
        is protected; 

    EECommonBlocks(me:out; 
    	    aM:IDMapOfPaveBlockIMapOfPaveBlock from BOPTools) 
    	is protected; 
     
    EFCommonBlocks(me:out;  
    	     aMapCB:IDMapOfPaveBlockIMapOfInteger from BOPTools) 
        is protected;  
	 
    EENewVertices (me:out;  
    	    aM:IndexedDataMapOfShapeInteger from BooleanOperations) 
    	is protected;  

    EENewVertices (me:out;  
    	    aV:Vertex from TopoDS;  
    	    aM:IndexedDataMapOfShapeInteger from BooleanOperations) 
    	is protected; 
     
    EFNewVertices (me:out; 
    	    aM:IndexedDataMapOfShapeInteger from BooleanOperations) 
    	is protected; 
     
    EFNewVertices (me:out; 
    	    aV:Vertex from TopoDS;  
    	    aM:IndexedDataMapOfShapeInteger from BooleanOperations) 
    	is protected;   
	 
    UpdateCommonBlocks(me:out) 
    	is protected;  
     
    UpdatePaveBlocks(me:out) 
    	is protected; 
	 
    SplitIndex(me; 
    	    aPB:PaveBlock from BOPTools) 
	returns Integer from Standard  
    	is protected;		     
    	 
    MakeBlocks(me:out) 
    	is protected;   

    -------------------------------------------------------------- 
    ---	  
    ---  Some API FUNCTIONS  
    ---  	    	 
    SplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  

    SplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	
    SplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	
    SplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	
    SplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	
    SplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
     
    SplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
     
    SplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
     
    SplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  

    SplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  
    --
    SplitsFace  (me:out;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools) 
    	returns Integer from Standard;  

    SplitsFace  (me:out;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  

    CommonBlocksFace (me:out;  
    	         nF  :Integer from Standard;  
    	         aLCB:out ListOfCommonBlock from NMTTools) 
    	returns Integer from Standard;   
	
    PrepareFace(me:out;  
    	    nF  :  Integer from Standard; 
    	    aF  : out Face from TopoDS); 
     
    -- 
    RealPaveBlock(me:out;   
    	    aPB:PaveBlock from BOPTools) 
	returns PaveBlock from BOPTools; 
    ---C++: return const & 	 
    -- 
    RealSplitsFace  (me:out;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
	 
    HasRealSplitsInOnFace (me:out; 
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard) 
    	returns Boolean from Standard; 
	 
    RealSplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
     
    RealSplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
     
    RealSplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
     
    RealSplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 

    RealSplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from BOPTools); 
    --   
    PrepareSetForFace(me:out;   
    	    	nF1 :Integer from Standard;  
    	        nF2 :Integer from Standard;
    	    	aPSF:out PaveSet from BOPTools); 
		 
    PutPaveOnCurve(me:out;   
    	    	aPSF: PaveSet from BOPTools; 
		aTol: Real from Standard;  
		aBC : out Curve from BOPTools); 
	 
    PutBoundPaveOnCurve (me:out; 
    	    	    aBC :out Curve from BOPTools;	 
     	    	    aFF :out SSInterference from BOPTools); 
    	
    PutBoundPaveOnCurve (me:out;  
    	    	    aP  : Pnt from  gp; 
		    aT  : Real from Standard; 			 
    	    	    aBC :out Curve from BOPTools;	 
     	    	    aFF :out SSInterference from BOPTools); 
    	
    FindPave            (me:out; 
		    aP  : Pnt from gp;  
    	    	    aTpV: Real from Standard;  
    	    	    aPS : PaveSet from BOPTools; 
		    aPV :out Pave from BOPTools) 
    	returns Boolean from Standard; 
	 
    CheckIntermediatePoint(me:out;  
    	    	    aPB : PaveBlock      from BOPTools;  
    	    	    aPBR: PaveBlock      from BOPTools;  
     	    	    aTol: Real  from  Standard) 
    	returns Integer from Standard; 	
		
    IsExistingPaveBlock (me:out; 
    	    	    aPB : PaveBlock      from BOPTools; 
     	    	    aFF : SSInterference from BOPTools) 
    	returns Boolean from Standard;  
	 
    MakePCurves (me:out); 
     
fields 
    myIntrPool         :  PInterferencePool from BOPTools    	is protected; 
    myDS               :  PShapesDataStructure from NMTDS   	is protected;   
    myIsDone           :  Boolean from Standard                 is protected; 
    myNbSources        :  Integer from Standard                 is protected;  
    myNbEdges          :  Integer from Standard           	is protected;      
    myDSIt             :  IteratorOfCoupleOfShape from NMTTools is protected;
    -- 
    myPavePool         :  PavePool from BOPTools                is protected;     
    myPavePoolNew      :  PavePool from BOPTools                is protected;  
    myCommonBlockPool  :  CommonBlockPool from NMTTools         is protected;  
    mySplitShapesPool  :  SplitShapesPool from BOPTools	        is protected;    
    -- 
    myContext          :  Context from IntTools                 is protected; 
    mySectionAttribute :  SSIntersectionAttribute from BOPTools is protected;
end PaveFiller;
