// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
//
-- File:	GEOMAlgo.cdl
-- Created:	Sat Dec 04 12:36:22 2004
-- Author:	Peter KURNEV
--		<peter@PREFEX>
---Copyright:	 Matra Datavision 2004


package GEOMAlgo 

	---Purpose: 

uses  
    TCollection, 
    TColStd, 
    Geom,     
    Bnd, 
    gp,	  
    GeomAdaptor,
    TopAbs,
    TopoDS, 
    TopTools, 
    IntTools, 
    BOPTools, 
    BOP     
    
is   
    --  enumerations 
    --
    enumeration State is 
    	ST_UNKNOWN, 
	ST_IN,
	ST_OUT,
	ST_ON, 
	ST_ONIN, 
	ST_ONOUT, 
	ST_INOUT    
    end State;
    -- 
    --  classes 
    -- 
    deferred class Algo;
    deferred class ShapeAlgo; 
    -- 
    --  gluer    	     
    class Gluer; 
    class GlueAnalyser; 
    class CoupleOfShapes; 
    class PassKey;  
    class PassKeyMapHasher; 
    class PassKeyShape;  
    class SurfaceTools; 
    class Tools;  
    
    --	     
    --  finder on 
    deferred class ShapeSolid;
    class WireSolid; 
    class ShellSolid; 
    class VertexSolid; 
    class SolidSolid; 
    class FinderShapeOn; 
    -- 
    class FinderShapeOn1;
    class StateCollector;
    --
    --  instantiations
    class IndexedDataMapOfPassKeyShapeListOfShape   
	instantiates IndexedDataMap from TCollection (PassKeyShape from GEOMAlgo, 
						      ListOfShape from TopTools, 
                                                      PassKeyMapHasher from GEOMAlgo); 
     
    class IndexedDataMapOfShapeBox  
    	instantiates IndexedDataMap from TCollection   	(Shape from TopoDS,
	    		    		         	 Box from Bnd,
	    		    		         	 ShapeMapHasher from TopTools);
    class IndexedDataMapOfIntegerShape  
    	instantiates IndexedDataMap from TCollection   	(Integer from Standard,
	    		    		         	 Shape from TopoDS,
	    		    		         	 MapIntegerHasher from TColStd); 
							  
    class ListOfCoupleOfShapes  
    	instantiates List from TCollection  (CoupleOfShapes from GEOMAlgo);


    class IndexedDataMapOfShapeState  
    	instantiates IndexedDataMap from TCollection   	(Shape from TopoDS,
	    		    		         	 State from TopAbs,  
	    	    	    	    	    	    	 ShapeMapHasher from TopTools);
--
    class ListOfPnt  
    	instantiates List from TCollection  (Pnt from gp);

--    class IndexedDataMapOfPassKeyInteger   
--	instantiates IndexedDataMap from TCollection (PassKeyRoot from GEOMAlgo, 
--						      Integer from Standard, 
--                                                      PassKeyMapHasher from GEOMAlgo); 
						       

    class DataMapOfPassKeyInteger   
	instantiates DataMap from TCollection (PassKey from GEOMAlgo, 
					       Integer from Standard, 
                                               PassKeyMapHasher from GEOMAlgo);


end GEOMAlgo;
