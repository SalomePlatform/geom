--  Copyright (C) 2007-2008  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
--  File:	NMTTools_CheckerSI.cdl
--  Created:	Mon Feb 19 11:23:55 2007
--  Author:	Peter KURNEV
--
class CheckerSI from NMTTools 
    	inherits PaveFiller from NMTTools 
	---Purpose: 

uses 
    ShapeEnum  from  TopAbs

--raises

is
 
    Create 
    	returns CheckerSI from NMTTools;  
    ---C++: alias "Standard_EXPORT virtual ~NMTTools_CheckerSI();" 
     
    Perform (me:out) 
	is redefined; 
	 
    Init  (me:out) 
    	is redefined protected;
 
    Clear (me:out) 
    	is redefined protected;
 
    PreparePaveBlocks (me:out;   
    	    nE:Integer from Standard) 
    	is redefined protected;  		

    PreparePaveBlocks (me:out; 
    	    aType1: ShapeEnum  from  TopAbs; 
    	    aType2: ShapeEnum  from  TopAbs) 
    	is redefined protected; 
    
    StopStatus(me) 
    	returns Integer from Standard;   


fields
    myStopStatus: Integer from Standard is protected; 
     
end CheckerSI;
