-- Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
-- 
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either 
-- version 2.1 of the License.
-- 
-- This library is distributed in the hope that it will be useful 
-- but WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public  
-- License along with this library; if not, write to the Free Software 
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
-- 
-- File:	NMTDS.cdl
-- Created:	Fri Nov 28 10:13:19 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>


package NMTDS 

	---Purpose: 

uses   
    
    TCollection, 
    TColStd,
    Bnd,
    TopoDS, 
    TopAbs, 
    TopTools, 
    BooleanOperations,
    BOPTColStd
is  
    class ShapesDataStructure;
    class IndexRange;   
    
    -- Modified to Add new classes Thu Sep 14 14:35:18 2006 
    -- Contribution of Samtech www.samcef.com BEGIN 
    class Iterator; 
    class PassKey; 
    class PassKeyBoolean; 
    class PassKeyMapHasher; 
    -- Contribution of Samtech www.samcef.com END  
    
    pointer PShapesDataStructure to ShapesDataStructure from NMTDS;

    class CArray1OfIndexRange instantiates 
	CArray1 from BOPTColStd(IndexRange from NMTDS); 
     
    class ListOfIndexedDataMapOfShapeAncestorsSuccessors instantiates 
	List from TCollection(IndexedDataMapOfShapeAncestorsSuccessors from BooleanOperations); 
	 
    class IndexedDataMapOfIntegerIndexedDataMapOfShapeInteger instantiates 
    	IndexedDataMap from TCollection(Integer        from Standard, 
	    	    	    	    	IndexedDataMapOfShapeInteger from BooleanOperations, 
					MapIntegerHasher from TColStd); 
    
    -- Modified to Add new classes Thu Sep 14 14:35:18 2006 
    -- Contribution of Samtech www.samcef.com BEGIN 
    class ListOfPassKey  instantiates 
	List from TCollection(PassKey from NMTDS);  
     
    class MapOfPassKey instantiates
    	Map from TCollection(PassKey from NMTDS, 
    	    	    	     PassKeyMapHasher from NMTDS);  
			     
    class ListOfPassKeyBoolean  instantiates 
	List from TCollection(PassKeyBoolean from NMTDS); 
     
    class MapOfPassKeyBoolean instantiates
    	Map from TCollection(PassKeyBoolean from NMTDS, 
    	    	    	     PassKeyMapHasher from NMTDS);   
    -- Contribution of Samtech www.samcef.com END


    class IndexedDataMapOfShapeBox  
    	instantiates IndexedDataMap from TCollection   	(Shape from TopoDS,
	    		    		         	 Box from Bnd,
	    		    		         	 ShapeMapHasher from TopTools);
    class IndexedDataMapOfIntegerShape  
    	instantiates IndexedDataMap from TCollection   	(Integer from Standard,
	    		    		         	 Shape from TopoDS,
	    		    		         	 MapIntegerHasher from TColStd); 

 
end NMTDS;
