// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
// See http://www.salome-platform.org/
//
-- File:	GEOMAlgo_CoupleOfShapes.cdl
-- Created:	Wed Dec 15 13:00:10 2004
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2004


class CoupleOfShapes from GEOMAlgo 

	---Purpose: 

uses
    Shape from TopoDS

--raises

is 
    Create 
    	returns CoupleOfShapes from GEOMAlgo; 

    SetShapes(me:out; 
    	    aS1: Shape from TopoDS; 
    	    aS2: Shape from TopoDS);
     
    SetShape1(me:out; 
    	    aS1: Shape from TopoDS); 
	 
    SetShape2(me:out; 
    	    aS2: Shape from TopoDS);     

    Shapes(me; 
    	    aS1:out Shape from TopoDS; 
    	    aS2:out Shape from TopoDS); 

    Shape1(me) 
    	returns Shape from TopoDS; 
    ---C++:return const &  
     
    Shape2(me) 
    	returns Shape from TopoDS; 
    ---C++:return const & 

fields  

    myShape1: Shape from TopoDS is protected;   
    myShape2: Shape from TopoDS is protected;   

end CoupleOfShapes;
