// Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
// CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Lesser General Public
// License as published by the Free Software Foundation; either 
// version 2.1 of the License.
// 
// This library is distributed in the hope that it will be useful 
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
// Lesser General Public License for more details.
//
// You should have received a copy of the GNU Lesser General Public  
// License along with this library; if not, write to the Free Software 
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
//
// See http://www.salome-platform.org/
//
-- File:	GEOMAlgo_WireSolid.cdl
-- Created:	Wed Jan 12 10:17:00 2005
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2005


class WireSolid from GEOMAlgo 
    	inherits ShapeSolid from GEOMAlgo
	---Purpose: 

--uses 
--raises

is 
    Create   
    	returns WireSolid from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_WireSolid();" 
    
    Perform (me:out) 
	is redefined; 
	 
    Prepare(me:out)  
   	 is redefined protected;
     
    BuildResult (me:out) 
	is redefined protected; 
    
--fields
    
end WireSolid;
