-- Copyright (C) 2007-2012  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	GEOMAlgo_WESCorrector.cdl
-- Created:	
-- Author:	Peter KURNEV
--
class WESCorrector from GEOMAlgo  
    inherits Algo from GEOMAlgo

	---Purpose: 
    	---  The algorithm to change the Wire Edges Set (WES) contents.
    	--   The NewWES will contain only wires instead of wires and edges. 
    	--
uses
    WireEdgeSet          from GEOMAlgo,
    PWireEdgeSet         from GEOMAlgo,
    ListOfConnexityBlock from BOP 
    
is 
    Create   
    	returns WESCorrector from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_WESCorrector();"  
    ---Purpose:  
    -- Empty constructor; 
    -- 
    
    SetWES  (me:out; 
		aWES: WireEdgeSet from GEOMAlgo);  
    ---Purpose: 
    -- Modifier 
    --
    Perform (me:out) 
    	is redefined; 
    ---Purpose: 
    --- Performs the algorithm that  consists  of  two  steps 
    --- 1. Make conexity blocks (  DoConnexityBlocks()  )     
    --- 2. Make corrections     (  DoCorrections()  )        
    ---
      
    WES     (me:out) 
    	returns WireEdgeSet from GEOMAlgo; 
    ---C++:  return &  
    ---Purpose: 
    --- Selector 
    ---
    NewWES  (me:out) 
    	returns WireEdgeSet from GEOMAlgo; 
    ---C++:  return &   
    ---Purpose: 
    --- Selector 
    ---
    DoConnexityBlocks(me:out) 
    	is protected; 
       
    DoCorrections(me:out) 
    	is protected; 

fields 

    myWES             : PWireEdgeSet         from GEOMAlgo is protected; 
    myNewWES          : WireEdgeSet          from GEOMAlgo is protected;  
    myConnexityBlocks : ListOfConnexityBlock from BOP is protected;  

end WESCorrector;
