--  Copyright (C) 2007-2008  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
-- 
-- File:	NMTDS_BndSphere.cdl
-- Created:	
-- Author:	Peter KURNEV
--		<pkv@irinox>


class BndSphere from NMTDS 

	---Purpose: 

uses
    Pnt from gp

is 
    Create 
    	returns BndSphere from NMTDS; 
    ---C++: alias "Standard_EXPORT virtual ~NMTDS_BndSphere();"  
     
    SetCenter(me:out; 
    	    theP:Pnt from gp); 
    ---C++: inline 
     
    Center(me) 
    	returns Pnt from gp; 
    ---C++:return const& 	
    ---C++: inline 
     
    SetRadius(me:out; 
    	    theR:Real from Standard);     
    ---C++: inline 
    
    Radius(me) 
    	returns Real from Standard; 
    ---C++: inline 
     
    SetGap(me:out; 
    	    theGap:Real from Standard);     
    ---C++: inline

    Gap(me) 
    	returns Real from Standard; 
    ---C++: inline

    Add(me:out;  
    	    theOther: BndSphere from NMTDS); 
    ---C++: inline	     

    IsOut(me;  
    	    theOther: BndSphere from NMTDS)  
    	returns Boolean from Standard;  

    SquareExtent(me)  
    	returns Real from Standard;
    ---C++: inline
fields 
    myCenter: Pnt from gp is protected;   
    myRadius: Real from Standard is protected;   
    myGap   : Real from Standard is protected;   

end BndSphere;
