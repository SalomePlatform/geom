-- File   :     Partition_Spliter.cdl
-- Created:     Thu Aug 02 16:07:39 2001
-- Author :     Benedicte MARTIN
---Copyright:    OPEN CASCADE  2001

class Spliter from Partition

        ---Purpose: Split solids, shells and  faces  into parts of the
        --          same  topology  if  reconstruction  level  is  not
        --          limited.

uses
    Inter3d             from Partition,
    Loop2d              from Partition,
    Builder             from BRep,
    ShapeEnum           from TopAbs,
    Compound            from TopoDS,
    Face                from TopoDS,
    Edge                from TopoDS,
    Shape               from TopoDS,
    MapOfOrientedShape  from TopTools,
    IndexedMapOfShape   from TopTools,
    DataMapOfShapeShape from TopTools,
    ListOfShape         from TopTools,
    MapOfShape          from TopTools,
    AsDes               from BRepAlgo,
    Image               from BRepAlgo

is
    Create  returns Spliter from Partition;
        ---Purpose: constructor

    AddShape ( me : in out; S : Shape from TopoDS);
        ---Purpose: add object Shape to be splitted.
        --          If S  is  a  COMPOUND  or  COMPSOLID,  it  will be
        --          exploded  in  order  to  get  more  simple  object
        --          shapes. 
        --          Object shapes that  are  vertices,  edges or wires
        --          won't be splitted and won't be in a result.

    AddTool  ( me : in out; S : Shape from TopoDS);
        ---Purpose: add cutting tool

    Compute (me : in out; Limit : ShapeEnum from TopAbs
                          = TopAbs_SHAPE);
        ---Purpose: produce a result which  is  a compound of parts of
        --          object shapes.  A  part  can  be  either a vertex,
        --          edge, wire, face, shell or solid.
        --          By default, a part is  of  the same topology as an
        --          object  shape,   else   <Limit>   restricts  parts
        --          reconstruction.
        --          If <Limit> == TopAbs_VERTEX, only new vertices are
        --          returned in the result

    KeepShapesInside (me : in out; S : Shape from TopoDS);
        ---Purpose: remove shapes that are outside of S from result.
        --          S should be an object shape.
        ---Warning: call it after Compute()

    RemoveShapesInside (me : in out; S : Shape from TopoDS);
        ---Purpose: remove shapes that are inside S from result.
        --          S should be an object shape.
        ---Warning: call it after Compute()

    Shape ( me ) returns Shape from TopoDS;
        ---Purpose: return resulting compound

    Clear ( me : in out);
        ---Purpose: clear fields


        ---Category: private methods


    MakeShells (me: in out; S : Shape from TopoDS;
                            NS: in out ListOfShape from TopTools) is private;
        ---Purpose: split S into shells

    MakeFaces (me: in out; S : Shape from TopoDS)
        returns Shape from TopoDS is private;
        ---Purpose: split faces of S, return compound of new faces

    MakeEdges (me; 
               E : Edge from TopoDS;
               VOnE : ListOfShape from TopTools;
               NE : in out ListOfShape from TopTools) 
        is private;
        ---Purpose: cut E by vertices  VOnE,  return list of new edges
        --          NE
    
    FindFacesInside (me: in out; S : Shape from TopoDS;
                                 CheckClosed : Boolean = Standard_False;
                                 All         : Boolean = Standard_False)
        returns Shape from TopoDS is private;
        ---Purpose: return compound of faces  of other shapes that are
        --          inside <S>. <S>  must  have image in myImageShape.
        --          <CheckClosed> makes avoid faces that do not form a
        --          closed shell
        --          <All> makes return already added faces

    CheckTool ( me: in out; S : Shape from TopoDS)
        returns Boolean from Standard is private;
        ---Purpose: Return True if <S>  is  a tool shape. Prepare tool
        --          faces of <S> for the search of internal faces.

    MergeEqualEdges (me: in out; LE : ListOfShape from TopTools) is private;
        ---Purpose: among LE, find  equal  edges,  choose ones to keep
        --          and make them have  pcurves  on all faces they are
        --          shared by
        --          <LE> contains edge splits

fields

    myDoneStep     : ShapeEnum           from TopAbs;   -- reconstructed topology
    myShape        : Compound            from TopoDS;   -- result
    myBuilder      : Builder             from BRep;
    		   			   
    myListShapes   : ListOfShape         from TopTools; -- object shapes
    myMapFaces     : MapOfShape          from TopTools; -- object faces
    myMapTools     : MapOfShape          from TopTools; -- tool faces
    myFaceShapeMap : DataMapOfShapeShape from TopTools; -- to find a shape by face
    		   			   
    myNewSection   : MapOfShape          from TopTools; -- new secton edges
		   			   
    myAsDes        : AsDes               from BRepAlgo;
    myImagesFaces  : Image               from BRepAlgo;   
    myImagesEdges  : Image               from BRepAlgo;    
    myImageShape   : Image               from BRepAlgo;
    
        -- contains info of same domain shapes and section edges
    myInter3d      : Inter3d             from Partition;
    
        -- avoid rebuilding twice commont part of solids
    myAddedFacesMap: MapOfOrientedShape  from TopTools;
    
        -- equal splits
    myEqualEdges   : MapOfShape          from TopTools;
    
        -- shape and its internal faces
    myInternalFaces: DataMapOfShapeShape from TopTools;
    
end Spliter;
