//  File      : GEOMDS_Application.cdl
//  Created   :
//  Author    : Yves FRICAUD
//  Project   : SALOME
//  Module    : GEOM
//  Copyright : OPEN CASCADE
//  $Header$


class Application from GEOMDS  inherits Application from TDocStd

	---Purpose: 

uses
    Label                    from TDF,
    SequenceOfExtendedString from TColStd,
    CString                  from Standard,
    Document                 from TDocStd


is

    Create 
    returns mutable Application from GEOMDS;
    
    Formats(me: mutable; Formats: out SequenceOfExtendedString from TColStd) 
    is redefined;    

    ResourcesName (me: mutable) returns CString from Standard;

end Application;
