-- Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
-- 
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either 
-- version 2.1 of the License.
-- 
-- This library is distributed in the hope that it will be useful 
-- but WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public  
-- License along with this library; if not, write to the Free Software 
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http:--www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
-- File:	GEOMAlgo_SolidSolid.cdl
-- Created:	Wed Jan 26 12:05:14 2005
-- Author:	Peter KURNEV
--		<pkv@irinox>
---Copyright:	 Matra Datavision 2005


class SolidSolid from GEOMAlgo 
    inherits ShellSolid from GEOMAlgo 
    
	---Purpose: 

uses 
    Shape from TopoDS

--raises

is
    Create   
    	returns SolidSolid from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_SolidSolid();" 
    
    Perform (me:out) 
	is redefined; 
	 
    BuildResult (me:out) 
	is redefined protected; 	
    
    SetShape2 (me:out;  
    	    aS: Shape from TopoDS);

    Shape2 (me)  
    	returns Shape from TopoDS; 
    ---C++: return const &  

fields
    myS2: Shape from TopoDS is protected; 
    
end SolidSolid;
