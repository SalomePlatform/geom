-- Copyright (C) 2005  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
-- 
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either 
-- version 2.1 of the License.
-- 
-- This library is distributed in the hope that it will be useful 
-- but WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public  
-- License along with this library; if not, write to the Free Software 
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http:--www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
-- File:	GEOMAlgo_Clsf.cdl
-- Created:	Wed Nov 22 10:19:29 2006
-- Author:	Peter KURNEV
--		<pkv@irinox>


deferred class Clsf from GEOMAlgo 
    inherits HAlgo from GEOMAlgo 
     
	---Purpose: 

uses 
    State from TopAbs,
    Pnt from gp, 
    Curve from Geom,
    Surface from Geom 
    
--raises

is 
    Initialize 
    	returns mutable Clsf from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_Clsf();"  
     
    SetPnt(me:mutable; 
    	    aP:Pnt from gp); 
	     
    Pnt(me) 
    	returns Pnt from gp; 
    ---C++:return const& 	 
	 
    SetTolerance(me:mutable; 
    	    aT:Real from Standard);  
	 
    Tolerance(me) 
    	returns Real from Standard;       
	 
    State(me) 
    	returns State from TopAbs; 
	 
    CanBeON(me; 
    	    aCT:Curve from Geom) 
	returns Boolean from Standard 
    	is virtual;     

    CanBeON(me; 
    	    aST:Surface from Geom) 
	returns Boolean from Standard 
    	is virtual;     
	
fields 
    myState    :State from TopAbs is protected;
    myPnt      :Pnt from gp is protected;
    myTolerance:Real from Standard is protected; 

end Clsf;
