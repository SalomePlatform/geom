--  Copyright (C) 2007-2011  CEA/DEN, EDF R&D, OPEN CASCADE
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2.1 of the License.
--
--  This library is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--  Lesser General Public License for more details.
--
--  You should have received a copy of the GNU Lesser General Public
--  License along with this library; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
--  See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--
-- File:	GEOMAlgo_WESScaler.cdl
-- Created:	
-- Author:	
--		<pkv@VORTEX>
 

class WESScaler from GEOMAlgo  
    	inherits Algo from GEOMAlgo  

	---Purpose: 

uses 
    Face from TopoDS, 
    Shape  from TopoDS,
    ListOfShape from  TopTools,	
    DataMapOfOrientedShapeShape from GEOMAlgo,
    WireEdgeSet from GEOMAlgo,  
    PWireEdgeSet from GEOMAlgo  
 
--raises

is 
    Create 
    	---Purpose: Empty constructor    
    	returns WESScaler from GEOMAlgo; 
    ---C++: alias "Standard_EXPORT virtual ~GEOMAlgo_WESScaler();"  
     
    SetScale  (me:out; 
		aWES: Real from Standard);  
    ---Purpose: 
    -- Modifier  
      
    Scale(me) 
	returns Real from Standard;       
    ---Purpose: 
    -- Selector  
    	 
    SetFace  (me:out; 
    	    	aF: Face from TopoDS); 
     
    Face (me) 
    	returns Face from TopoDS; 
    ---C++:  return const & 
     
    SetEdges  (me:out; 
		aLE:ListOfShape from  TopTools);  
     
    Edges  (me)
	 returns ListOfShape from  TopTools;  
    ---C++:  return const &		 
    
    Perform(me:out)  
    	---Purpose:  Performs the algorithm 
    	is redefined;   
      
    FaceScaled (me) 
    	returns Face from TopoDS; 
    ---C++:  return const & 
     
    EdgesScaled  (me)
	 returns ListOfShape from  TopTools;  
    ---C++:  return const &   
    
    Image(me; 
    	    aS:Shape from TopoDS)  
    	returns Shape from TopoDS; 
    ---C++: return const &  
    ---Purpose: 
     
    Origin(me; 
    	    aS:Shape from TopoDS)  
    	returns Shape from TopoDS; 
    ---C++: return const &   
    
    ---Purpose: 
    Images(me)  
    	returns  DataMapOfOrientedShapeShape from GEOMAlgo; 
    ---C++: return const &  
    ---Purpose: 
    --- Selector 
     
    Origins(me)  
    	returns   DataMapOfOrientedShapeShape from GEOMAlgo; 
    ---C++: return const &  
    ---Purpose: 
    --- Selector    
     
    CheckData(me:out)  
    	---Purpose:  Performs the algorithm 
    	is redefined protected; 
	 
fields 
    myScale         : Real from Standard is protected; 
    myFace          : Face from TopoDS is protected;    
    
    myEdges         : ListOfShape from  TopTools is protected;    
    myFaceScaled    : Face from TopoDS is protected;    
    myEdgesScaled   : ListOfShape from  TopTools is protected;
    myImages        : DataMapOfOrientedShapeShape from GEOMAlgo is protected;     
    myOrigins       : DataMapOfOrientedShapeShape from GEOMAlgo is protected;      
    myShapeTmp      : Shape  from TopoDS is protected;    
end WESScaler;

